module instr_fetch(pc, instruction, next_pc);

	input [15:0] pc;
	output [15:0] next_pc;
	output [15:0] instruction;



endmodule
