module instr_fetch(pc, instruction, new_pc);

	input [15:0] pc;
	output [15:0] new_pc;
	output [15:0] instruction;



endmodule
