library verilog;
use verilog.vl_types.all;
entity not1 is
    port(
        in1             : in     vl_logic;
        \out\           : out    vl_logic
    );
end not1;
