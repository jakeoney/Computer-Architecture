
module dff_207 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_206 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_189 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_190 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_191 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_192 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_193 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_194 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_195 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_196 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_197 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_198 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_199 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_200 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_201 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_173 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_174 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_175 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_176 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_177 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_178 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_179 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_180 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_181 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_182 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_183 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_184 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_185 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_186 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_187 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_188 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_157 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_158 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_159 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_160 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_161 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_162 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_163 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_164 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_165 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_166 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_167 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_168 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_169 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_170 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_171 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_172 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_205 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_204 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_203 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_202 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_156 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_155 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_154 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_153 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_152 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_151 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_150 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_149 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_148 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_147 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_146 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_145 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_144 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_143 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_142 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_141 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_140 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_139 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_138 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_137 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_136 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_135 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_134 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_133 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_132 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_131 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_130 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_129 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_128 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_127 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_126 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_125 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_124 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_123 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_122 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_121 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_120 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_119 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_118 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_117 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_116 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_115 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_114 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_113 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_112 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_111 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_110 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_109 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_108 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_107 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_106 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_105 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_104 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_103 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_102 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_101 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_100 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_99 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_98 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_97 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_96 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_95 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_94 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_93 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_92 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_91 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_90 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_89 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_88 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_87 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_86 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_85 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_84 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_83 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_82 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_81 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_80 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_79 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_78 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_77 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_76 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_75 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_74 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_73 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_72 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_71 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_70 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_69 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_68 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_67 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_66 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_65 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_64 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_63 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_62 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_61 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_60 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_59 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_58 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_57 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_56 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_55 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_54 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_53 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_52 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_51 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_50 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_49 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_48 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_47 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_46 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_45 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_44 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_43 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_42 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_41 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_40 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_39 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_38 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_37 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_36 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_35 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_34 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_33 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_32 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_31 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_30 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_29 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_28 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_27 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_26 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_25 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_24 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_23 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_22 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_21 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_20 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_19 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_18 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_17 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_16 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_15 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_14 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_13 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_12 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_11 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_10 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_9 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_8 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_7 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_6 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_5 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_4 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_0 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_1 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_2 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_3 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module memc_Size16_3 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, n214, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n1162), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n1161), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n1160), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n1159), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n1158), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n1157), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n1156), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n1155), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n1154), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1153), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1152), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1151), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1150), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1149), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1148), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1147), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n1146), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n1145), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n1144), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n1143), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n1142), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n1141), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n1140), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n1139), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1138), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1137), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1136), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1135), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1134), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1133), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1132), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1131), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n1130), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n1129), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n1128), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n1127), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n1126), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n1125), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n1124), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n1123), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1122), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1121), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1120), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1119), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1118), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1117), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1116), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1115), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n1114), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n1113), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n1112), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n1111), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n1110), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n1109), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n1108), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n1107), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1106), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1105), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1104), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1103), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1102), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1101), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1100), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1099), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n1098), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n1097), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n1096), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n1095), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n1094), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n1093), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n1092), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n1091), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1090), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1089), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1088), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1087), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1086), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1085), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1084), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1083), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n1082), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n1081), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n1080), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n1079), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n1078), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n1077), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n1076), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n1075), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1074), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1073), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1072), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1071), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1070), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1069), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1068), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1067), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n1066), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n1065), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n1064), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n1063), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n1062), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n1061), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n1060), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n1059), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1058), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1057), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1056), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1055), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1054), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1053), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1052), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1051), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n1050), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n1049), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n1048), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n1047), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n1046), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n1045), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n1044), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n1043), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1042), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1041), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1040), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1039), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1038), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1037), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1036), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1035), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n1034), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n1033), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n1032), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n1031), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n1030), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n1029), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n1028), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n1027), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1026), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1025), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1024), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1023), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1022), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1021), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1020), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1019), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n1018), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n1017), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n1016), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n1015), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n1014), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n1013), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n1012), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n1011), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n1010), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n1009), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n1008), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n1007), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n1006), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n1005), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n1004), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n1003), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n1002), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n1001), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n1000), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n999), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n998), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n997), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n996), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n995), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n994), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n993), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n992), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n991), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n990), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n989), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n988), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n987), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n986), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n985), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n984), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n983), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n982), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n981), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n980), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n979), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n978), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n977), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n976), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n975), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n974), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n973), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n972), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n971), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n970), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n969), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n968), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n967), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n966), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n965), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n964), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n963), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n962), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n961), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n960), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n959), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n958), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n957), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n956), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n955), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n954), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n953), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n952), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n951), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n950), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n949), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n948), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n947), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n946), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n945), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n944), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n943), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n942), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n941), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n940), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n939), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n938), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n937), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n936), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n935), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n934), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n933), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n932), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n931), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n930), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n929), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n928), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n927), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n926), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n925), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n924), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n923), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n922), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n921), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n920), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n919), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n918), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n917), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n916), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n915), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n914), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n913), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n912), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n911), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n910), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n909), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n908), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n907), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n906), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n905), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n904), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n903), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n902), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n901), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n900), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n899), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n898), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n897), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n896), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n895), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n894), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n893), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n892), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n891), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n890), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n889), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n888), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n887), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n886), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n885), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n884), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n883), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n882), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n881), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n880), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n879), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n878), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n877), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n876), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n875), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n874), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n873), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n872), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n871), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n870), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n869), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n868), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n867), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n866), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n865), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n864), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n863), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n862), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n861), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n860), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n859), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n858), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n857), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n856), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n855), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n854), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n853), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n852), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n851), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n850), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n849), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n848), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n847), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n846), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n845), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n844), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n843), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n842), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n841), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n840), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n839), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n838), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n837), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n836), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n835), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n834), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n833), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n832), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n831), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n830), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n829), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n828), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n827), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n826), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n825), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n824), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n823), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n822), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n821), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n820), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n819), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n818), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n817), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n816), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n815), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n814), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n813), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n812), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n811), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n810), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n809), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n808), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n807), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n806), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n805), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n804), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n803), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n802), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n801), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n800), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n799), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n798), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n797), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n796), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n795), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n794), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n793), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n792), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n791), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n790), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n789), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n788), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n787), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n786), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n785), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n784), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n783), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n782), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n781), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n780), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n779), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n778), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n777), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n776), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n775), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n774), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n773), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n772), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n771), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n770), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n769), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n768), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n767), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n766), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n765), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n764), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n763), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n762), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n761), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n760), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n759), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n758), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n757), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n756), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n755), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n754), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n753), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n752), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n751), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n750), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n749), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n748), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n747), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n746), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n745), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n744), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n743), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n742), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n741), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n740), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n739), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n738), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n737), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n736), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n735), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n734), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n733), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n732), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n731), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n730), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n729), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n728), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n727), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n726), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n725), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n724), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n723), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n722), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n721), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n720), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n719), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n718), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n717), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n716), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n715), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n714), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n713), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n712), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n711), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n710), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n709), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n708), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n707), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n706), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n705), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n704), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n703), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n702), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n701), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n700), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n699), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n698), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n697), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n696), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n695), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n694), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n693), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n692), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n691), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n690), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n689), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n688), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n687), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n686), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n685), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n684), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n683), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n682), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n681), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n680), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n679), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n678), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n677), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n676), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n675), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n674), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n673), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n672), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n671), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n670), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n669), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n668), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n667), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n666), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n665), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n664), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n663), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n662), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n661), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n660), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n659), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n658), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n657), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n656), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n655), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n654), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n653), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n652), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n651), .CLK(clk), .Q(\mem<31><0> ) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n214) );
  INVX2 U2 ( .A(n1225), .Y(n1207) );
  INVX1 U3 ( .A(n1209), .Y(n1217) );
  INVX1 U4 ( .A(n1208), .Y(n1214) );
  INVX1 U5 ( .A(n1209), .Y(n1215) );
  INVX1 U6 ( .A(n1208), .Y(n1221) );
  INVX1 U7 ( .A(n1208), .Y(n1220) );
  INVX1 U8 ( .A(n1208), .Y(n1210) );
  INVX1 U9 ( .A(n1207), .Y(n1212) );
  INVX1 U10 ( .A(n1208), .Y(n1219) );
  INVX1 U11 ( .A(n1209), .Y(n1216) );
  INVX4 U12 ( .A(n44), .Y(n45) );
  INVX4 U13 ( .A(n42), .Y(n43) );
  INVX4 U14 ( .A(n40), .Y(n41) );
  INVX4 U15 ( .A(n38), .Y(n39) );
  INVX4 U16 ( .A(n36), .Y(n37) );
  INVX4 U17 ( .A(n34), .Y(n35) );
  INVX4 U18 ( .A(n32), .Y(n33) );
  INVX4 U19 ( .A(n30), .Y(n31) );
  INVX4 U20 ( .A(n28), .Y(n29) );
  INVX4 U21 ( .A(n26), .Y(n27) );
  INVX4 U22 ( .A(n24), .Y(n25) );
  INVX4 U23 ( .A(n22), .Y(n23) );
  INVX1 U24 ( .A(n1169), .Y(N32) );
  INVX1 U25 ( .A(n1170), .Y(N31) );
  INVX1 U26 ( .A(n1172), .Y(N29) );
  INVX1 U27 ( .A(n1173), .Y(N28) );
  INVX1 U28 ( .A(n1174), .Y(N27) );
  INVX1 U29 ( .A(n1175), .Y(N26) );
  INVX1 U30 ( .A(n1176), .Y(N25) );
  INVX1 U31 ( .A(n1177), .Y(N24) );
  INVX1 U32 ( .A(n1178), .Y(N23) );
  INVX1 U33 ( .A(n1179), .Y(N22) );
  INVX1 U34 ( .A(n1180), .Y(N21) );
  INVX1 U35 ( .A(n1181), .Y(N20) );
  INVX1 U36 ( .A(n1182), .Y(N19) );
  INVX1 U37 ( .A(n1183), .Y(N18) );
  INVX1 U38 ( .A(n1184), .Y(N17) );
  INVX1 U39 ( .A(n1308), .Y(n1224) );
  INVX1 U40 ( .A(n1308), .Y(n1225) );
  INVX1 U41 ( .A(n1225), .Y(n1209) );
  INVX1 U42 ( .A(n1224), .Y(n1208) );
  INVX1 U43 ( .A(n1195), .Y(n1196) );
  INVX1 U44 ( .A(n1195), .Y(n1197) );
  INVX2 U45 ( .A(n1207), .Y(n1213) );
  INVX1 U46 ( .A(n1195), .Y(n1198) );
  INVX1 U47 ( .A(n1195), .Y(n1199) );
  INVX2 U48 ( .A(n1195), .Y(n1200) );
  INVX2 U49 ( .A(n1207), .Y(n1218) );
  INVX2 U50 ( .A(n1195), .Y(n1201) );
  INVX1 U51 ( .A(n1188), .Y(n1191) );
  INVX1 U52 ( .A(n1194), .Y(n1202) );
  INVX2 U53 ( .A(n1207), .Y(n1222) );
  INVX1 U54 ( .A(n1194), .Y(n1203) );
  INVX1 U55 ( .A(n1194), .Y(n1204) );
  INVX1 U56 ( .A(n1194), .Y(n1205) );
  INVX2 U57 ( .A(n1194), .Y(n1206) );
  INVX1 U58 ( .A(n1188), .Y(n1193) );
  INVX1 U59 ( .A(n1171), .Y(N30) );
  INVX1 U60 ( .A(n1309), .Y(n1195) );
  INVX1 U61 ( .A(N14), .Y(n1315) );
  INVX1 U62 ( .A(n1311), .Y(n1188) );
  INVX2 U63 ( .A(n1207), .Y(n1211) );
  INVX2 U64 ( .A(n1207), .Y(n1223) );
  INVX1 U65 ( .A(n1312), .Y(n1190) );
  INVX1 U66 ( .A(n1188), .Y(n1189) );
  INVX1 U67 ( .A(n1188), .Y(n1192) );
  INVX1 U68 ( .A(n1313), .Y(n1186) );
  INVX1 U69 ( .A(n1313), .Y(n1187) );
  INVX8 U70 ( .A(n1273), .Y(n1272) );
  INVX1 U71 ( .A(n1315), .Y(n1185) );
  INVX1 U72 ( .A(n1309), .Y(n1194) );
  INVX1 U73 ( .A(n117), .Y(n1253) );
  INVX1 U74 ( .A(n119), .Y(n1269) );
  INVX1 U75 ( .A(n118), .Y(n1254) );
  INVX1 U76 ( .A(n116), .Y(n1242) );
  INVX1 U77 ( .A(rst), .Y(n1307) );
  INVX4 U78 ( .A(n60), .Y(n102) );
  BUFX2 U79 ( .A(n101), .Y(n1) );
  BUFX2 U80 ( .A(n99), .Y(n2) );
  BUFX2 U81 ( .A(n97), .Y(n3) );
  BUFX2 U82 ( .A(n95), .Y(n4) );
  BUFX2 U83 ( .A(n91), .Y(n5) );
  BUFX2 U84 ( .A(n89), .Y(n6) );
  BUFX2 U85 ( .A(n87), .Y(n7) );
  BUFX2 U86 ( .A(n85), .Y(n8) );
  BUFX2 U87 ( .A(n83), .Y(n9) );
  BUFX2 U88 ( .A(n81), .Y(n10) );
  BUFX2 U89 ( .A(n64), .Y(n11) );
  BUFX2 U90 ( .A(n93), .Y(n12) );
  BUFX2 U91 ( .A(n59), .Y(n13) );
  BUFX2 U92 ( .A(n57), .Y(n14) );
  BUFX2 U93 ( .A(n55), .Y(n15) );
  BUFX2 U94 ( .A(n53), .Y(n16) );
  BUFX2 U95 ( .A(n51), .Y(n17) );
  BUFX2 U96 ( .A(n49), .Y(n18) );
  BUFX2 U97 ( .A(n47), .Y(n19) );
  INVX4 U98 ( .A(n1274), .Y(n1270) );
  INVX2 U99 ( .A(n1316), .Y(n20) );
  INVX2 U100 ( .A(n1316), .Y(n21) );
  INVX1 U101 ( .A(n1316), .Y(n1317) );
  INVX1 U102 ( .A(N13), .Y(n1313) );
  AND2X2 U103 ( .A(n1271), .B(n142), .Y(n22) );
  AND2X2 U104 ( .A(n1271), .B(n144), .Y(n24) );
  AND2X2 U105 ( .A(n1271), .B(n146), .Y(n26) );
  AND2X2 U106 ( .A(n1271), .B(n117), .Y(n28) );
  AND2X2 U107 ( .A(n1271), .B(n148), .Y(n30) );
  AND2X2 U108 ( .A(n1271), .B(n150), .Y(n32) );
  AND2X2 U109 ( .A(n1271), .B(n152), .Y(n34) );
  AND2X2 U110 ( .A(n1271), .B(n154), .Y(n36) );
  AND2X2 U111 ( .A(n1271), .B(n156), .Y(n38) );
  AND2X2 U112 ( .A(n1271), .B(n158), .Y(n40) );
  AND2X2 U113 ( .A(n1271), .B(n160), .Y(n42) );
  AND2X2 U114 ( .A(n1271), .B(n119), .Y(n44) );
  AND2X2 U115 ( .A(n1271), .B(n162), .Y(n46) );
  INVX1 U116 ( .A(n46), .Y(n47) );
  AND2X2 U117 ( .A(n1271), .B(n164), .Y(n48) );
  INVX1 U118 ( .A(n48), .Y(n49) );
  AND2X2 U119 ( .A(n1271), .B(n166), .Y(n50) );
  INVX1 U120 ( .A(n50), .Y(n51) );
  AND2X2 U121 ( .A(n1271), .B(n168), .Y(n52) );
  INVX1 U122 ( .A(n52), .Y(n53) );
  AND2X2 U123 ( .A(n1271), .B(n170), .Y(n54) );
  INVX1 U124 ( .A(n54), .Y(n55) );
  AND2X2 U125 ( .A(n1271), .B(n172), .Y(n56) );
  INVX1 U126 ( .A(n56), .Y(n57) );
  AND2X2 U127 ( .A(n1271), .B(n174), .Y(n58) );
  INVX1 U128 ( .A(n58), .Y(n59) );
  AND2X2 U129 ( .A(n1272), .B(n118), .Y(n60) );
  AND2X2 U130 ( .A(n1307), .B(n1227), .Y(n61) );
  AND2X2 U131 ( .A(\data_in<0> ), .B(n1272), .Y(n62) );
  AND2X2 U132 ( .A(n1270), .B(n120), .Y(n63) );
  INVX1 U133 ( .A(n63), .Y(n64) );
  AND2X2 U134 ( .A(\data_in<1> ), .B(n1272), .Y(n65) );
  AND2X2 U135 ( .A(\data_in<2> ), .B(n1272), .Y(n66) );
  AND2X2 U136 ( .A(\data_in<3> ), .B(n1272), .Y(n67) );
  AND2X2 U137 ( .A(\data_in<4> ), .B(n1272), .Y(n68) );
  AND2X2 U138 ( .A(\data_in<5> ), .B(n1272), .Y(n69) );
  AND2X2 U139 ( .A(\data_in<6> ), .B(n1272), .Y(n70) );
  AND2X2 U140 ( .A(\data_in<7> ), .B(n1272), .Y(n71) );
  AND2X2 U141 ( .A(\data_in<8> ), .B(n1272), .Y(n72) );
  AND2X2 U142 ( .A(\data_in<9> ), .B(n1272), .Y(n73) );
  AND2X2 U143 ( .A(\data_in<10> ), .B(n1272), .Y(n74) );
  AND2X2 U144 ( .A(\data_in<11> ), .B(n1272), .Y(n75) );
  AND2X2 U145 ( .A(\data_in<12> ), .B(n1272), .Y(n76) );
  AND2X2 U146 ( .A(\data_in<13> ), .B(n1272), .Y(n77) );
  AND2X2 U147 ( .A(\data_in<14> ), .B(n1272), .Y(n78) );
  AND2X2 U148 ( .A(\data_in<15> ), .B(n1272), .Y(n79) );
  AND2X2 U149 ( .A(n1270), .B(n122), .Y(n80) );
  INVX1 U150 ( .A(n80), .Y(n81) );
  AND2X2 U151 ( .A(n1270), .B(n124), .Y(n82) );
  INVX1 U152 ( .A(n82), .Y(n83) );
  AND2X2 U153 ( .A(n1270), .B(n126), .Y(n84) );
  INVX1 U154 ( .A(n84), .Y(n85) );
  AND2X2 U155 ( .A(n1270), .B(n128), .Y(n86) );
  INVX1 U156 ( .A(n86), .Y(n87) );
  AND2X2 U157 ( .A(n1270), .B(n130), .Y(n88) );
  INVX1 U158 ( .A(n88), .Y(n89) );
  AND2X2 U159 ( .A(n1270), .B(n132), .Y(n90) );
  INVX1 U160 ( .A(n90), .Y(n91) );
  AND2X2 U161 ( .A(n1270), .B(n116), .Y(n92) );
  INVX1 U162 ( .A(n92), .Y(n93) );
  AND2X2 U163 ( .A(n1270), .B(n134), .Y(n94) );
  INVX1 U164 ( .A(n94), .Y(n95) );
  AND2X2 U165 ( .A(n1270), .B(n136), .Y(n96) );
  INVX1 U166 ( .A(n96), .Y(n97) );
  AND2X2 U167 ( .A(n1270), .B(n138), .Y(n98) );
  INVX1 U168 ( .A(n98), .Y(n99) );
  AND2X2 U169 ( .A(n1270), .B(n140), .Y(n100) );
  INVX1 U170 ( .A(n100), .Y(n101) );
  INVX1 U171 ( .A(n61), .Y(n1274) );
  INVX4 U172 ( .A(n61), .Y(n1273) );
  INVX1 U173 ( .A(n1310), .Y(n1309) );
  AND2X1 U174 ( .A(n1311), .B(n1309), .Y(n103) );
  INVX1 U175 ( .A(n1312), .Y(n1311) );
  AND2X1 U176 ( .A(n214), .B(n1314), .Y(n104) );
  INVX1 U177 ( .A(n1315), .Y(n1314) );
  BUFX2 U178 ( .A(n64), .Y(n1228) );
  BUFX2 U179 ( .A(n64), .Y(n1229) );
  BUFX2 U180 ( .A(n81), .Y(n1230) );
  BUFX2 U181 ( .A(n81), .Y(n1231) );
  BUFX2 U182 ( .A(n83), .Y(n1232) );
  BUFX2 U183 ( .A(n83), .Y(n1233) );
  BUFX2 U184 ( .A(n85), .Y(n1234) );
  BUFX2 U185 ( .A(n85), .Y(n1235) );
  BUFX2 U186 ( .A(n87), .Y(n1236) );
  BUFX2 U187 ( .A(n87), .Y(n1237) );
  BUFX2 U188 ( .A(n89), .Y(n1238) );
  BUFX2 U189 ( .A(n89), .Y(n1239) );
  BUFX2 U190 ( .A(n91), .Y(n1240) );
  BUFX2 U191 ( .A(n91), .Y(n1241) );
  BUFX2 U192 ( .A(n93), .Y(n1243) );
  BUFX2 U193 ( .A(n93), .Y(n1244) );
  BUFX2 U194 ( .A(n95), .Y(n1245) );
  BUFX2 U195 ( .A(n95), .Y(n1246) );
  BUFX2 U196 ( .A(n97), .Y(n1247) );
  BUFX2 U197 ( .A(n97), .Y(n1248) );
  BUFX2 U198 ( .A(n99), .Y(n1249) );
  BUFX2 U199 ( .A(n99), .Y(n1250) );
  BUFX2 U200 ( .A(n101), .Y(n1251) );
  BUFX2 U201 ( .A(n101), .Y(n1252) );
  BUFX2 U202 ( .A(n1350), .Y(n105) );
  INVX1 U203 ( .A(n105), .Y(n1742) );
  BUFX2 U204 ( .A(n1367), .Y(n106) );
  INVX1 U205 ( .A(n106), .Y(n1759) );
  BUFX2 U206 ( .A(n1384), .Y(n107) );
  INVX1 U207 ( .A(n107), .Y(n1776) );
  BUFX2 U208 ( .A(n1401), .Y(n108) );
  INVX1 U209 ( .A(n108), .Y(n1793) );
  BUFX2 U210 ( .A(n1418), .Y(n109) );
  INVX1 U211 ( .A(n109), .Y(n1810) );
  BUFX2 U212 ( .A(n1579), .Y(n110) );
  INVX1 U213 ( .A(n110), .Y(n1692) );
  BUFX2 U214 ( .A(n1709), .Y(n111) );
  INVX1 U215 ( .A(n111), .Y(n1827) );
  AND2X1 U216 ( .A(n1216), .B(n103), .Y(n112) );
  AND2X1 U217 ( .A(n1187), .B(n104), .Y(n113) );
  AND2X1 U218 ( .A(n1308), .B(n103), .Y(n114) );
  AND2X1 U219 ( .A(n1313), .B(n104), .Y(n115) );
  AND2X1 U220 ( .A(n113), .B(n1828), .Y(n116) );
  AND2X1 U221 ( .A(n1828), .B(n115), .Y(n117) );
  AND2X1 U222 ( .A(n1828), .B(n1692), .Y(n118) );
  AND2X1 U223 ( .A(n1828), .B(n1827), .Y(n119) );
  AND2X1 U224 ( .A(n112), .B(n113), .Y(n120) );
  INVX1 U225 ( .A(n120), .Y(n121) );
  AND2X1 U226 ( .A(n113), .B(n114), .Y(n122) );
  INVX1 U227 ( .A(n122), .Y(n123) );
  AND2X1 U228 ( .A(n113), .B(n1742), .Y(n124) );
  INVX1 U229 ( .A(n124), .Y(n125) );
  AND2X1 U230 ( .A(n113), .B(n1759), .Y(n126) );
  INVX1 U231 ( .A(n126), .Y(n127) );
  AND2X1 U232 ( .A(n113), .B(n1776), .Y(n128) );
  INVX1 U233 ( .A(n128), .Y(n129) );
  AND2X1 U234 ( .A(n113), .B(n1793), .Y(n130) );
  INVX1 U235 ( .A(n130), .Y(n131) );
  AND2X1 U236 ( .A(n113), .B(n1810), .Y(n132) );
  INVX1 U237 ( .A(n132), .Y(n133) );
  AND2X1 U238 ( .A(n112), .B(n115), .Y(n134) );
  INVX1 U239 ( .A(n134), .Y(n135) );
  AND2X1 U240 ( .A(n114), .B(n115), .Y(n136) );
  INVX1 U241 ( .A(n136), .Y(n137) );
  AND2X1 U242 ( .A(n1742), .B(n115), .Y(n138) );
  INVX1 U243 ( .A(n138), .Y(n139) );
  AND2X1 U244 ( .A(n1759), .B(n115), .Y(n140) );
  INVX1 U245 ( .A(n140), .Y(n141) );
  AND2X1 U246 ( .A(n1776), .B(n115), .Y(n142) );
  INVX1 U247 ( .A(n142), .Y(n143) );
  AND2X1 U248 ( .A(n1793), .B(n115), .Y(n144) );
  INVX1 U249 ( .A(n144), .Y(n145) );
  AND2X1 U250 ( .A(n1810), .B(n115), .Y(n146) );
  INVX1 U251 ( .A(n146), .Y(n147) );
  AND2X1 U252 ( .A(n112), .B(n1692), .Y(n148) );
  INVX1 U253 ( .A(n148), .Y(n149) );
  AND2X1 U254 ( .A(n114), .B(n1692), .Y(n150) );
  INVX1 U255 ( .A(n150), .Y(n151) );
  AND2X1 U256 ( .A(n1742), .B(n1692), .Y(n152) );
  INVX1 U257 ( .A(n152), .Y(n153) );
  AND2X1 U258 ( .A(n1759), .B(n1692), .Y(n154) );
  INVX1 U259 ( .A(n154), .Y(n155) );
  AND2X1 U260 ( .A(n1776), .B(n1692), .Y(n156) );
  INVX1 U261 ( .A(n156), .Y(n157) );
  AND2X1 U262 ( .A(n1793), .B(n1692), .Y(n158) );
  INVX1 U263 ( .A(n158), .Y(n159) );
  AND2X1 U264 ( .A(n1810), .B(n1692), .Y(n160) );
  INVX1 U265 ( .A(n160), .Y(n161) );
  AND2X1 U266 ( .A(n112), .B(n1827), .Y(n162) );
  INVX1 U267 ( .A(n162), .Y(n163) );
  BUFX2 U268 ( .A(n47), .Y(n1255) );
  BUFX2 U269 ( .A(n47), .Y(n1256) );
  AND2X1 U270 ( .A(n114), .B(n1827), .Y(n164) );
  INVX1 U271 ( .A(n164), .Y(n165) );
  BUFX2 U272 ( .A(n49), .Y(n1257) );
  BUFX2 U273 ( .A(n49), .Y(n1258) );
  AND2X1 U274 ( .A(n1742), .B(n1827), .Y(n166) );
  INVX1 U275 ( .A(n166), .Y(n167) );
  BUFX2 U276 ( .A(n51), .Y(n1259) );
  BUFX2 U277 ( .A(n51), .Y(n1260) );
  AND2X1 U278 ( .A(n1759), .B(n1827), .Y(n168) );
  INVX1 U279 ( .A(n168), .Y(n169) );
  BUFX2 U280 ( .A(n53), .Y(n1261) );
  BUFX2 U281 ( .A(n53), .Y(n1262) );
  AND2X1 U282 ( .A(n1776), .B(n1827), .Y(n170) );
  INVX1 U283 ( .A(n170), .Y(n171) );
  BUFX2 U284 ( .A(n55), .Y(n1263) );
  BUFX2 U285 ( .A(n55), .Y(n1264) );
  AND2X1 U286 ( .A(n1793), .B(n1827), .Y(n172) );
  INVX1 U287 ( .A(n172), .Y(n173) );
  BUFX2 U288 ( .A(n57), .Y(n1265) );
  BUFX2 U289 ( .A(n57), .Y(n1266) );
  AND2X1 U290 ( .A(n1810), .B(n1827), .Y(n174) );
  INVX1 U291 ( .A(n174), .Y(n175) );
  BUFX2 U292 ( .A(n59), .Y(n1267) );
  BUFX2 U293 ( .A(n59), .Y(n1268) );
  MUX2X1 U294 ( .B(n177), .A(n178), .S(n1196), .Y(n176) );
  MUX2X1 U295 ( .B(n180), .A(n181), .S(n1196), .Y(n179) );
  MUX2X1 U296 ( .B(n183), .A(n184), .S(n1196), .Y(n182) );
  MUX2X1 U297 ( .B(n186), .A(n187), .S(n1196), .Y(n185) );
  MUX2X1 U298 ( .B(n189), .A(n190), .S(n1187), .Y(n188) );
  MUX2X1 U299 ( .B(n192), .A(n193), .S(n1196), .Y(n191) );
  MUX2X1 U300 ( .B(n195), .A(n196), .S(n1196), .Y(n194) );
  MUX2X1 U301 ( .B(n198), .A(n199), .S(n1196), .Y(n197) );
  MUX2X1 U302 ( .B(n201), .A(n202), .S(n1196), .Y(n200) );
  MUX2X1 U303 ( .B(n204), .A(n205), .S(n1187), .Y(n203) );
  MUX2X1 U304 ( .B(n207), .A(n208), .S(n1197), .Y(n206) );
  MUX2X1 U305 ( .B(n210), .A(n211), .S(n1197), .Y(n209) );
  MUX2X1 U306 ( .B(n213), .A(n215), .S(n1197), .Y(n212) );
  MUX2X1 U307 ( .B(n217), .A(n218), .S(n1197), .Y(n216) );
  MUX2X1 U308 ( .B(n220), .A(n221), .S(n1187), .Y(n219) );
  MUX2X1 U309 ( .B(n223), .A(n224), .S(n1197), .Y(n222) );
  MUX2X1 U310 ( .B(n226), .A(n227), .S(n1197), .Y(n225) );
  MUX2X1 U311 ( .B(n229), .A(n230), .S(n1197), .Y(n228) );
  MUX2X1 U312 ( .B(n232), .A(n233), .S(n1197), .Y(n231) );
  MUX2X1 U313 ( .B(n235), .A(n236), .S(n1187), .Y(n234) );
  MUX2X1 U314 ( .B(n238), .A(n239), .S(n1197), .Y(n237) );
  MUX2X1 U315 ( .B(n241), .A(n242), .S(n1197), .Y(n240) );
  MUX2X1 U316 ( .B(n244), .A(n245), .S(n1197), .Y(n243) );
  MUX2X1 U317 ( .B(n247), .A(n248), .S(n1197), .Y(n246) );
  MUX2X1 U318 ( .B(n250), .A(n251), .S(n1187), .Y(n249) );
  MUX2X1 U319 ( .B(n253), .A(n254), .S(n1198), .Y(n252) );
  MUX2X1 U320 ( .B(n256), .A(n257), .S(n1198), .Y(n255) );
  MUX2X1 U321 ( .B(n259), .A(n260), .S(n1198), .Y(n258) );
  MUX2X1 U322 ( .B(n262), .A(n263), .S(n1198), .Y(n261) );
  MUX2X1 U323 ( .B(n265), .A(n266), .S(n1187), .Y(n264) );
  MUX2X1 U324 ( .B(n268), .A(n269), .S(n1198), .Y(n267) );
  MUX2X1 U325 ( .B(n271), .A(n272), .S(n1198), .Y(n270) );
  MUX2X1 U326 ( .B(n274), .A(n275), .S(n1198), .Y(n273) );
  MUX2X1 U327 ( .B(n277), .A(n278), .S(n1198), .Y(n276) );
  MUX2X1 U328 ( .B(n280), .A(n281), .S(n1187), .Y(n279) );
  MUX2X1 U329 ( .B(n283), .A(n284), .S(n1198), .Y(n282) );
  MUX2X1 U330 ( .B(n286), .A(n287), .S(n1198), .Y(n285) );
  MUX2X1 U331 ( .B(n289), .A(n290), .S(n1198), .Y(n288) );
  MUX2X1 U332 ( .B(n292), .A(n293), .S(n1198), .Y(n291) );
  MUX2X1 U333 ( .B(n295), .A(n296), .S(n1187), .Y(n294) );
  MUX2X1 U334 ( .B(n298), .A(n299), .S(n1199), .Y(n297) );
  MUX2X1 U335 ( .B(n301), .A(n302), .S(n1199), .Y(n300) );
  MUX2X1 U336 ( .B(n304), .A(n305), .S(n1199), .Y(n303) );
  MUX2X1 U337 ( .B(n307), .A(n308), .S(n1199), .Y(n306) );
  MUX2X1 U338 ( .B(n310), .A(n311), .S(n1187), .Y(n309) );
  MUX2X1 U339 ( .B(n313), .A(n314), .S(n1199), .Y(n312) );
  MUX2X1 U340 ( .B(n316), .A(n317), .S(n1199), .Y(n315) );
  MUX2X1 U341 ( .B(n319), .A(n320), .S(n1199), .Y(n318) );
  MUX2X1 U342 ( .B(n322), .A(n323), .S(n1199), .Y(n321) );
  MUX2X1 U343 ( .B(n325), .A(n326), .S(n1187), .Y(n324) );
  MUX2X1 U344 ( .B(n328), .A(n329), .S(n1199), .Y(n327) );
  MUX2X1 U345 ( .B(n331), .A(n332), .S(n1199), .Y(n330) );
  MUX2X1 U346 ( .B(n334), .A(n335), .S(n1199), .Y(n333) );
  MUX2X1 U347 ( .B(n337), .A(n338), .S(n1199), .Y(n336) );
  MUX2X1 U348 ( .B(n340), .A(n341), .S(n1187), .Y(n339) );
  MUX2X1 U349 ( .B(n343), .A(n344), .S(n1200), .Y(n342) );
  MUX2X1 U350 ( .B(n346), .A(n347), .S(n1200), .Y(n345) );
  MUX2X1 U351 ( .B(n349), .A(n350), .S(n1200), .Y(n348) );
  MUX2X1 U352 ( .B(n352), .A(n353), .S(n1200), .Y(n351) );
  MUX2X1 U353 ( .B(n355), .A(n356), .S(n1187), .Y(n354) );
  MUX2X1 U354 ( .B(n358), .A(n359), .S(n1200), .Y(n357) );
  MUX2X1 U355 ( .B(n361), .A(n362), .S(n1200), .Y(n360) );
  MUX2X1 U356 ( .B(n364), .A(n365), .S(n1200), .Y(n363) );
  MUX2X1 U357 ( .B(n367), .A(n368), .S(n1200), .Y(n366) );
  MUX2X1 U358 ( .B(n370), .A(n371), .S(n1186), .Y(n369) );
  MUX2X1 U359 ( .B(n373), .A(n374), .S(n1200), .Y(n372) );
  MUX2X1 U360 ( .B(n376), .A(n377), .S(n1200), .Y(n375) );
  MUX2X1 U361 ( .B(n379), .A(n380), .S(n1200), .Y(n378) );
  MUX2X1 U362 ( .B(n382), .A(n383), .S(n1200), .Y(n381) );
  MUX2X1 U363 ( .B(n385), .A(n386), .S(n1186), .Y(n384) );
  MUX2X1 U364 ( .B(n388), .A(n389), .S(n1201), .Y(n387) );
  MUX2X1 U365 ( .B(n391), .A(n392), .S(n1201), .Y(n390) );
  MUX2X1 U366 ( .B(n394), .A(n395), .S(n1201), .Y(n393) );
  MUX2X1 U367 ( .B(n397), .A(n398), .S(n1201), .Y(n396) );
  MUX2X1 U368 ( .B(n400), .A(n401), .S(n1186), .Y(n399) );
  MUX2X1 U369 ( .B(n403), .A(n404), .S(n1201), .Y(n402) );
  MUX2X1 U370 ( .B(n406), .A(n407), .S(n1201), .Y(n405) );
  MUX2X1 U371 ( .B(n409), .A(n410), .S(n1201), .Y(n408) );
  MUX2X1 U372 ( .B(n412), .A(n413), .S(n1201), .Y(n411) );
  MUX2X1 U373 ( .B(n415), .A(n416), .S(n1186), .Y(n414) );
  MUX2X1 U374 ( .B(n418), .A(n419), .S(n1201), .Y(n417) );
  MUX2X1 U375 ( .B(n421), .A(n422), .S(n1201), .Y(n420) );
  MUX2X1 U376 ( .B(n424), .A(n425), .S(n1201), .Y(n423) );
  MUX2X1 U377 ( .B(n427), .A(n428), .S(n1201), .Y(n426) );
  MUX2X1 U378 ( .B(n430), .A(n431), .S(n1186), .Y(n429) );
  MUX2X1 U379 ( .B(n433), .A(n434), .S(n1202), .Y(n432) );
  MUX2X1 U380 ( .B(n436), .A(n437), .S(n1202), .Y(n435) );
  MUX2X1 U381 ( .B(n439), .A(n440), .S(n1202), .Y(n438) );
  MUX2X1 U382 ( .B(n442), .A(n443), .S(n1202), .Y(n441) );
  MUX2X1 U383 ( .B(n445), .A(n446), .S(n1186), .Y(n444) );
  MUX2X1 U384 ( .B(n448), .A(n449), .S(n1202), .Y(n447) );
  MUX2X1 U385 ( .B(n451), .A(n452), .S(n1202), .Y(n450) );
  MUX2X1 U386 ( .B(n454), .A(n455), .S(n1202), .Y(n453) );
  MUX2X1 U387 ( .B(n457), .A(n458), .S(n1202), .Y(n456) );
  MUX2X1 U388 ( .B(n460), .A(n461), .S(n1186), .Y(n459) );
  MUX2X1 U389 ( .B(n463), .A(n464), .S(n1202), .Y(n462) );
  MUX2X1 U390 ( .B(n466), .A(n467), .S(n1202), .Y(n465) );
  MUX2X1 U391 ( .B(n469), .A(n470), .S(n1202), .Y(n468) );
  MUX2X1 U392 ( .B(n472), .A(n473), .S(n1202), .Y(n471) );
  MUX2X1 U393 ( .B(n475), .A(n476), .S(n1186), .Y(n474) );
  MUX2X1 U394 ( .B(n478), .A(n479), .S(n1203), .Y(n477) );
  MUX2X1 U395 ( .B(n481), .A(n482), .S(n1203), .Y(n480) );
  MUX2X1 U396 ( .B(n484), .A(n485), .S(n1203), .Y(n483) );
  MUX2X1 U397 ( .B(n487), .A(n488), .S(n1203), .Y(n486) );
  MUX2X1 U398 ( .B(n490), .A(n491), .S(n1186), .Y(n489) );
  MUX2X1 U399 ( .B(n493), .A(n494), .S(n1203), .Y(n492) );
  MUX2X1 U400 ( .B(n496), .A(n497), .S(n1203), .Y(n495) );
  MUX2X1 U401 ( .B(n499), .A(n500), .S(n1203), .Y(n498) );
  MUX2X1 U402 ( .B(n502), .A(n503), .S(n1203), .Y(n501) );
  MUX2X1 U403 ( .B(n505), .A(n506), .S(n1186), .Y(n504) );
  MUX2X1 U404 ( .B(n508), .A(n509), .S(n1203), .Y(n507) );
  MUX2X1 U405 ( .B(n511), .A(n512), .S(n1203), .Y(n510) );
  MUX2X1 U406 ( .B(n514), .A(n515), .S(n1203), .Y(n513) );
  MUX2X1 U407 ( .B(n517), .A(n518), .S(n1203), .Y(n516) );
  MUX2X1 U408 ( .B(n520), .A(n521), .S(n1186), .Y(n519) );
  MUX2X1 U409 ( .B(n523), .A(n524), .S(n1204), .Y(n522) );
  MUX2X1 U410 ( .B(n526), .A(n527), .S(n1204), .Y(n525) );
  MUX2X1 U411 ( .B(n529), .A(n530), .S(n1204), .Y(n528) );
  MUX2X1 U412 ( .B(n532), .A(n533), .S(n1204), .Y(n531) );
  MUX2X1 U413 ( .B(n535), .A(n536), .S(n1186), .Y(n534) );
  MUX2X1 U414 ( .B(n538), .A(n539), .S(n1204), .Y(n537) );
  MUX2X1 U415 ( .B(n541), .A(n542), .S(n1204), .Y(n540) );
  MUX2X1 U416 ( .B(n544), .A(n545), .S(n1204), .Y(n543) );
  MUX2X1 U417 ( .B(n547), .A(n548), .S(n1204), .Y(n546) );
  MUX2X1 U418 ( .B(n550), .A(n551), .S(n1187), .Y(n549) );
  MUX2X1 U419 ( .B(n553), .A(n554), .S(n1204), .Y(n552) );
  MUX2X1 U420 ( .B(n556), .A(n557), .S(n1204), .Y(n555) );
  MUX2X1 U421 ( .B(n559), .A(n560), .S(n1204), .Y(n558) );
  MUX2X1 U422 ( .B(n562), .A(n563), .S(n1204), .Y(n561) );
  MUX2X1 U423 ( .B(n565), .A(n566), .S(n1186), .Y(n564) );
  MUX2X1 U424 ( .B(n568), .A(n569), .S(n1205), .Y(n567) );
  MUX2X1 U425 ( .B(n571), .A(n572), .S(n1205), .Y(n570) );
  MUX2X1 U426 ( .B(n574), .A(n575), .S(n1205), .Y(n573) );
  MUX2X1 U427 ( .B(n577), .A(n578), .S(n1205), .Y(n576) );
  MUX2X1 U428 ( .B(n580), .A(n581), .S(n1187), .Y(n579) );
  MUX2X1 U429 ( .B(n583), .A(n584), .S(n1205), .Y(n582) );
  MUX2X1 U430 ( .B(n586), .A(n587), .S(n1205), .Y(n585) );
  MUX2X1 U431 ( .B(n589), .A(n590), .S(n1205), .Y(n588) );
  MUX2X1 U432 ( .B(n592), .A(n593), .S(n1205), .Y(n591) );
  MUX2X1 U433 ( .B(n595), .A(n596), .S(n1186), .Y(n594) );
  MUX2X1 U434 ( .B(n598), .A(n599), .S(n1205), .Y(n597) );
  MUX2X1 U435 ( .B(n601), .A(n602), .S(n1205), .Y(n600) );
  MUX2X1 U436 ( .B(n604), .A(n605), .S(n1205), .Y(n603) );
  MUX2X1 U437 ( .B(n607), .A(n608), .S(n1205), .Y(n606) );
  MUX2X1 U438 ( .B(n610), .A(n611), .S(n1186), .Y(n609) );
  MUX2X1 U439 ( .B(n613), .A(n614), .S(n1206), .Y(n612) );
  MUX2X1 U440 ( .B(n616), .A(n617), .S(n1206), .Y(n615) );
  MUX2X1 U441 ( .B(n619), .A(n620), .S(n1206), .Y(n618) );
  MUX2X1 U442 ( .B(n622), .A(n623), .S(n1206), .Y(n621) );
  MUX2X1 U443 ( .B(n625), .A(n626), .S(n1186), .Y(n624) );
  MUX2X1 U444 ( .B(n628), .A(n629), .S(n1206), .Y(n627) );
  MUX2X1 U445 ( .B(n631), .A(n632), .S(n1206), .Y(n630) );
  MUX2X1 U446 ( .B(n634), .A(n635), .S(n1206), .Y(n633) );
  MUX2X1 U447 ( .B(n637), .A(n638), .S(n1206), .Y(n636) );
  MUX2X1 U448 ( .B(n640), .A(n641), .S(n1186), .Y(n639) );
  MUX2X1 U449 ( .B(n643), .A(n644), .S(n1206), .Y(n642) );
  MUX2X1 U450 ( .B(n646), .A(n647), .S(n1206), .Y(n645) );
  MUX2X1 U451 ( .B(n649), .A(n650), .S(n1206), .Y(n648) );
  MUX2X1 U452 ( .B(n1164), .A(n1165), .S(n1206), .Y(n1163) );
  MUX2X1 U453 ( .B(n1167), .A(n1168), .S(n1186), .Y(n1166) );
  MUX2X1 U454 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n1211), .Y(n178) );
  MUX2X1 U455 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n1223), .Y(n177) );
  MUX2X1 U456 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n1211), .Y(n181) );
  MUX2X1 U457 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n1222), .Y(n180) );
  MUX2X1 U458 ( .B(n179), .A(n176), .S(n1193), .Y(n190) );
  MUX2X1 U459 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n1210), .Y(n184) );
  MUX2X1 U460 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n1210), .Y(n183) );
  MUX2X1 U461 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n1210), .Y(n187) );
  MUX2X1 U462 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n1210), .Y(n186) );
  MUX2X1 U463 ( .B(n185), .A(n182), .S(n1193), .Y(n189) );
  MUX2X1 U464 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n1210), .Y(n193) );
  MUX2X1 U465 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n1210), .Y(n192) );
  MUX2X1 U466 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n1210), .Y(n196) );
  MUX2X1 U467 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n1210), .Y(n195) );
  MUX2X1 U468 ( .B(n194), .A(n191), .S(n1193), .Y(n205) );
  MUX2X1 U469 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n1210), .Y(n199) );
  MUX2X1 U470 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n1210), .Y(n198) );
  MUX2X1 U471 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n1210), .Y(n202) );
  MUX2X1 U472 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n1210), .Y(n201) );
  MUX2X1 U473 ( .B(n200), .A(n197), .S(n1193), .Y(n204) );
  MUX2X1 U474 ( .B(n203), .A(n188), .S(n1185), .Y(n1169) );
  MUX2X1 U475 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n1211), .Y(n208) );
  MUX2X1 U476 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n1211), .Y(n207) );
  MUX2X1 U477 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n1211), .Y(n211) );
  MUX2X1 U478 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n1211), .Y(n210) );
  MUX2X1 U479 ( .B(n209), .A(n206), .S(n1193), .Y(n221) );
  MUX2X1 U480 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n1211), .Y(n215) );
  MUX2X1 U481 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n1211), .Y(n213) );
  MUX2X1 U482 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n1211), .Y(n218) );
  MUX2X1 U483 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n1211), .Y(n217) );
  MUX2X1 U484 ( .B(n216), .A(n212), .S(n1193), .Y(n220) );
  MUX2X1 U485 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n1211), .Y(n224) );
  MUX2X1 U486 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n1211), .Y(n223) );
  MUX2X1 U487 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n1211), .Y(n227) );
  MUX2X1 U488 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n1211), .Y(n226) );
  MUX2X1 U489 ( .B(n225), .A(n222), .S(n1193), .Y(n236) );
  MUX2X1 U490 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n1212), .Y(n230) );
  MUX2X1 U491 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n1212), .Y(n229) );
  MUX2X1 U492 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n1212), .Y(n233) );
  MUX2X1 U493 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n1212), .Y(n232) );
  MUX2X1 U494 ( .B(n231), .A(n228), .S(n1193), .Y(n235) );
  MUX2X1 U495 ( .B(n234), .A(n219), .S(n1185), .Y(n1170) );
  MUX2X1 U496 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n1212), .Y(n239) );
  MUX2X1 U497 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n1212), .Y(n238) );
  MUX2X1 U498 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n1212), .Y(n242) );
  MUX2X1 U499 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n1212), .Y(n241) );
  MUX2X1 U500 ( .B(n240), .A(n237), .S(n1193), .Y(n251) );
  MUX2X1 U501 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n1212), .Y(n245) );
  MUX2X1 U502 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n1212), .Y(n244) );
  MUX2X1 U503 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n1212), .Y(n248) );
  MUX2X1 U504 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n1212), .Y(n247) );
  MUX2X1 U505 ( .B(n246), .A(n243), .S(n1193), .Y(n250) );
  MUX2X1 U506 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n1213), .Y(n254) );
  MUX2X1 U507 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n1213), .Y(n253) );
  MUX2X1 U508 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n1213), .Y(n257) );
  MUX2X1 U509 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n1213), .Y(n256) );
  MUX2X1 U510 ( .B(n255), .A(n252), .S(n1193), .Y(n266) );
  MUX2X1 U511 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n1213), .Y(n260) );
  MUX2X1 U512 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n1213), .Y(n259) );
  MUX2X1 U513 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n1213), .Y(n263) );
  MUX2X1 U514 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n1213), .Y(n262) );
  MUX2X1 U515 ( .B(n261), .A(n258), .S(n1193), .Y(n265) );
  MUX2X1 U516 ( .B(n264), .A(n249), .S(n1185), .Y(n1171) );
  MUX2X1 U517 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n1213), .Y(n269) );
  MUX2X1 U518 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n1213), .Y(n268) );
  MUX2X1 U519 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n1213), .Y(n272) );
  MUX2X1 U520 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n1213), .Y(n271) );
  MUX2X1 U521 ( .B(n270), .A(n267), .S(n1192), .Y(n281) );
  MUX2X1 U522 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n1214), .Y(n275) );
  MUX2X1 U523 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n1214), .Y(n274) );
  MUX2X1 U524 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n1214), .Y(n278) );
  MUX2X1 U525 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n1214), .Y(n277) );
  MUX2X1 U526 ( .B(n276), .A(n273), .S(n1192), .Y(n280) );
  MUX2X1 U527 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n1214), .Y(n284) );
  MUX2X1 U528 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n1214), .Y(n283) );
  MUX2X1 U529 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n1214), .Y(n287) );
  MUX2X1 U530 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n1214), .Y(n286) );
  MUX2X1 U531 ( .B(n285), .A(n282), .S(n1192), .Y(n296) );
  MUX2X1 U532 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n1214), .Y(n290) );
  MUX2X1 U533 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n1214), .Y(n289) );
  MUX2X1 U534 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n1214), .Y(n293) );
  MUX2X1 U535 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n1214), .Y(n292) );
  MUX2X1 U536 ( .B(n291), .A(n288), .S(n1192), .Y(n295) );
  MUX2X1 U537 ( .B(n294), .A(n279), .S(n1185), .Y(n1172) );
  MUX2X1 U538 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n1215), .Y(n299) );
  MUX2X1 U539 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n1215), .Y(n298) );
  MUX2X1 U540 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n1215), .Y(n302) );
  MUX2X1 U541 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n1215), .Y(n301) );
  MUX2X1 U542 ( .B(n300), .A(n297), .S(n1192), .Y(n311) );
  MUX2X1 U543 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n1215), .Y(n305) );
  MUX2X1 U544 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n1215), .Y(n304) );
  MUX2X1 U545 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n1215), .Y(n308) );
  MUX2X1 U546 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n1215), .Y(n307) );
  MUX2X1 U547 ( .B(n306), .A(n303), .S(n1192), .Y(n310) );
  MUX2X1 U548 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n1215), .Y(n314) );
  MUX2X1 U549 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n1215), .Y(n313) );
  MUX2X1 U550 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n1215), .Y(n317) );
  MUX2X1 U551 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n1215), .Y(n316) );
  MUX2X1 U552 ( .B(n315), .A(n312), .S(n1192), .Y(n326) );
  MUX2X1 U553 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n1216), .Y(n320) );
  MUX2X1 U554 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n1216), .Y(n319) );
  MUX2X1 U555 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n1216), .Y(n323) );
  MUX2X1 U556 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n1216), .Y(n322) );
  MUX2X1 U557 ( .B(n321), .A(n318), .S(n1192), .Y(n325) );
  MUX2X1 U558 ( .B(n324), .A(n309), .S(n1185), .Y(n1173) );
  MUX2X1 U559 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n1216), .Y(n329) );
  MUX2X1 U560 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n1216), .Y(n328) );
  MUX2X1 U561 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n1216), .Y(n332) );
  MUX2X1 U562 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n1216), .Y(n331) );
  MUX2X1 U563 ( .B(n330), .A(n327), .S(n1192), .Y(n341) );
  MUX2X1 U564 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n1216), .Y(n335) );
  MUX2X1 U565 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n1216), .Y(n334) );
  MUX2X1 U566 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n1216), .Y(n338) );
  MUX2X1 U567 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n1216), .Y(n337) );
  MUX2X1 U568 ( .B(n336), .A(n333), .S(n1192), .Y(n340) );
  MUX2X1 U569 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n1217), .Y(n344) );
  MUX2X1 U570 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n1217), .Y(n343) );
  MUX2X1 U571 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n1217), .Y(n347) );
  MUX2X1 U572 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n1217), .Y(n346) );
  MUX2X1 U573 ( .B(n345), .A(n342), .S(n1192), .Y(n356) );
  MUX2X1 U574 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n1217), .Y(n350) );
  MUX2X1 U575 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n1217), .Y(n349) );
  MUX2X1 U576 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n1217), .Y(n353) );
  MUX2X1 U577 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n1217), .Y(n352) );
  MUX2X1 U578 ( .B(n351), .A(n348), .S(n1192), .Y(n355) );
  MUX2X1 U579 ( .B(n354), .A(n339), .S(n1185), .Y(n1174) );
  MUX2X1 U580 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n1217), .Y(n359) );
  MUX2X1 U581 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n1217), .Y(n358) );
  MUX2X1 U582 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n1217), .Y(n362) );
  MUX2X1 U583 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n1217), .Y(n361) );
  MUX2X1 U584 ( .B(n360), .A(n357), .S(n1191), .Y(n371) );
  MUX2X1 U585 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n1221), .Y(n365) );
  MUX2X1 U586 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n1220), .Y(n364) );
  MUX2X1 U587 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n1219), .Y(n368) );
  MUX2X1 U588 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n1218), .Y(n367) );
  MUX2X1 U589 ( .B(n366), .A(n363), .S(n1191), .Y(n370) );
  MUX2X1 U590 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n1222), .Y(n374) );
  MUX2X1 U591 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n1211), .Y(n373) );
  MUX2X1 U592 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n1211), .Y(n377) );
  MUX2X1 U593 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n1214), .Y(n376) );
  MUX2X1 U594 ( .B(n375), .A(n372), .S(n1191), .Y(n386) );
  MUX2X1 U595 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n1213), .Y(n380) );
  MUX2X1 U596 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n1210), .Y(n379) );
  MUX2X1 U597 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n1217), .Y(n383) );
  MUX2X1 U598 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n1215), .Y(n382) );
  MUX2X1 U599 ( .B(n381), .A(n378), .S(n1191), .Y(n385) );
  MUX2X1 U600 ( .B(n384), .A(n369), .S(n1185), .Y(n1175) );
  MUX2X1 U601 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n1218), .Y(n389) );
  MUX2X1 U602 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n1218), .Y(n388) );
  MUX2X1 U603 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n1218), .Y(n392) );
  MUX2X1 U604 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n1218), .Y(n391) );
  MUX2X1 U605 ( .B(n390), .A(n387), .S(n1191), .Y(n401) );
  MUX2X1 U606 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n1218), .Y(n395) );
  MUX2X1 U607 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n1218), .Y(n394) );
  MUX2X1 U608 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n1218), .Y(n398) );
  MUX2X1 U609 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n1218), .Y(n397) );
  MUX2X1 U610 ( .B(n396), .A(n393), .S(n1191), .Y(n400) );
  MUX2X1 U611 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n1218), .Y(n404) );
  MUX2X1 U612 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n1218), .Y(n403) );
  MUX2X1 U613 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n1218), .Y(n407) );
  MUX2X1 U614 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n1218), .Y(n406) );
  MUX2X1 U615 ( .B(n405), .A(n402), .S(n1191), .Y(n416) );
  MUX2X1 U616 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n1219), .Y(n410) );
  MUX2X1 U617 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n1219), .Y(n409) );
  MUX2X1 U618 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n1219), .Y(n413) );
  MUX2X1 U619 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n1219), .Y(n412) );
  MUX2X1 U620 ( .B(n411), .A(n408), .S(n1191), .Y(n415) );
  MUX2X1 U621 ( .B(n414), .A(n399), .S(n1185), .Y(n1176) );
  MUX2X1 U622 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n1219), .Y(n419) );
  MUX2X1 U623 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n1219), .Y(n418) );
  MUX2X1 U624 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n1219), .Y(n422) );
  MUX2X1 U625 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n1219), .Y(n421) );
  MUX2X1 U626 ( .B(n420), .A(n417), .S(n1191), .Y(n431) );
  MUX2X1 U627 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n1219), .Y(n425) );
  MUX2X1 U628 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n1219), .Y(n424) );
  MUX2X1 U629 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n1219), .Y(n428) );
  MUX2X1 U630 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n1219), .Y(n427) );
  MUX2X1 U631 ( .B(n426), .A(n423), .S(n1191), .Y(n430) );
  MUX2X1 U632 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n1220), .Y(n434) );
  MUX2X1 U633 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n1220), .Y(n433) );
  MUX2X1 U634 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n1220), .Y(n437) );
  MUX2X1 U635 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n1220), .Y(n436) );
  MUX2X1 U636 ( .B(n435), .A(n432), .S(n1191), .Y(n446) );
  MUX2X1 U637 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n1220), .Y(n440) );
  MUX2X1 U638 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n1220), .Y(n439) );
  MUX2X1 U639 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n1220), .Y(n443) );
  MUX2X1 U640 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n1220), .Y(n442) );
  MUX2X1 U641 ( .B(n441), .A(n438), .S(n1191), .Y(n445) );
  MUX2X1 U642 ( .B(n444), .A(n429), .S(n1185), .Y(n1177) );
  MUX2X1 U643 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n1220), .Y(n449) );
  MUX2X1 U644 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n1220), .Y(n448) );
  MUX2X1 U645 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n1220), .Y(n452) );
  MUX2X1 U646 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n1220), .Y(n451) );
  MUX2X1 U647 ( .B(n450), .A(n447), .S(n1190), .Y(n461) );
  MUX2X1 U648 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n1221), .Y(n455) );
  MUX2X1 U649 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n1221), .Y(n454) );
  MUX2X1 U650 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n1221), .Y(n458) );
  MUX2X1 U651 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n1221), .Y(n457) );
  MUX2X1 U652 ( .B(n456), .A(n453), .S(n1190), .Y(n460) );
  MUX2X1 U653 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n1221), .Y(n464) );
  MUX2X1 U654 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n1221), .Y(n463) );
  MUX2X1 U655 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n1221), .Y(n467) );
  MUX2X1 U656 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n1221), .Y(n466) );
  MUX2X1 U657 ( .B(n465), .A(n462), .S(n1190), .Y(n476) );
  MUX2X1 U658 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n1221), .Y(n470) );
  MUX2X1 U659 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n1221), .Y(n469) );
  MUX2X1 U660 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n1221), .Y(n473) );
  MUX2X1 U661 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n1221), .Y(n472) );
  MUX2X1 U662 ( .B(n471), .A(n468), .S(n1190), .Y(n475) );
  MUX2X1 U663 ( .B(n474), .A(n459), .S(n1185), .Y(n1178) );
  MUX2X1 U664 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n1222), .Y(n479) );
  MUX2X1 U665 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n1222), .Y(n478) );
  MUX2X1 U666 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n1222), .Y(n482) );
  MUX2X1 U667 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n1222), .Y(n481) );
  MUX2X1 U668 ( .B(n480), .A(n477), .S(n1190), .Y(n491) );
  MUX2X1 U669 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n1222), .Y(n485) );
  MUX2X1 U670 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n1222), .Y(n484) );
  MUX2X1 U671 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n1222), .Y(n488) );
  MUX2X1 U672 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n1222), .Y(n487) );
  MUX2X1 U673 ( .B(n486), .A(n483), .S(n1190), .Y(n490) );
  MUX2X1 U674 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n1222), .Y(n494) );
  MUX2X1 U675 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n1222), .Y(n493) );
  MUX2X1 U676 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n1222), .Y(n497) );
  MUX2X1 U677 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n1222), .Y(n496) );
  MUX2X1 U678 ( .B(n495), .A(n492), .S(n1190), .Y(n506) );
  MUX2X1 U679 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n1213), .Y(n500) );
  MUX2X1 U680 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n1222), .Y(n499) );
  MUX2X1 U681 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n1213), .Y(n503) );
  MUX2X1 U682 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n1217), .Y(n502) );
  MUX2X1 U683 ( .B(n501), .A(n498), .S(n1190), .Y(n505) );
  MUX2X1 U684 ( .B(n504), .A(n489), .S(n1185), .Y(n1179) );
  MUX2X1 U685 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n1217), .Y(n509) );
  MUX2X1 U686 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n1211), .Y(n508) );
  MUX2X1 U687 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n1211), .Y(n512) );
  MUX2X1 U688 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n1215), .Y(n511) );
  MUX2X1 U689 ( .B(n510), .A(n507), .S(n1190), .Y(n521) );
  MUX2X1 U690 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n1214), .Y(n515) );
  MUX2X1 U691 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n1215), .Y(n514) );
  MUX2X1 U692 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n1214), .Y(n518) );
  MUX2X1 U693 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n1220), .Y(n517) );
  MUX2X1 U694 ( .B(n516), .A(n513), .S(n1190), .Y(n520) );
  MUX2X1 U695 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n1222), .Y(n524) );
  MUX2X1 U696 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n1213), .Y(n523) );
  MUX2X1 U697 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n1222), .Y(n527) );
  MUX2X1 U698 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n1213), .Y(n526) );
  MUX2X1 U699 ( .B(n525), .A(n522), .S(n1190), .Y(n536) );
  MUX2X1 U700 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n1211), .Y(n530) );
  MUX2X1 U701 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n1211), .Y(n529) );
  MUX2X1 U702 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n1213), .Y(n533) );
  MUX2X1 U703 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n1211), .Y(n532) );
  MUX2X1 U704 ( .B(n531), .A(n528), .S(n1190), .Y(n535) );
  MUX2X1 U705 ( .B(n534), .A(n519), .S(n1185), .Y(n1180) );
  MUX2X1 U706 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n1211), .Y(n539) );
  MUX2X1 U707 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n1223), .Y(n538) );
  MUX2X1 U708 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n1213), .Y(n542) );
  MUX2X1 U709 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n1213), .Y(n541) );
  MUX2X1 U710 ( .B(n540), .A(n537), .S(n1189), .Y(n551) );
  MUX2X1 U711 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n1218), .Y(n545) );
  MUX2X1 U712 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n1223), .Y(n544) );
  MUX2X1 U713 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n1218), .Y(n548) );
  MUX2X1 U714 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n1213), .Y(n547) );
  MUX2X1 U715 ( .B(n546), .A(n543), .S(n1189), .Y(n550) );
  MUX2X1 U716 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n1223), .Y(n554) );
  MUX2X1 U717 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n1218), .Y(n553) );
  MUX2X1 U718 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n1222), .Y(n557) );
  MUX2X1 U719 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n1223), .Y(n556) );
  MUX2X1 U720 ( .B(n555), .A(n552), .S(n1189), .Y(n566) );
  MUX2X1 U721 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n1223), .Y(n560) );
  MUX2X1 U722 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n1213), .Y(n559) );
  MUX2X1 U723 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n1218), .Y(n563) );
  MUX2X1 U724 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n1211), .Y(n562) );
  MUX2X1 U725 ( .B(n561), .A(n558), .S(n1189), .Y(n565) );
  MUX2X1 U726 ( .B(n564), .A(n549), .S(n1185), .Y(n1181) );
  MUX2X1 U727 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n1211), .Y(n569) );
  MUX2X1 U728 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n1223), .Y(n568) );
  MUX2X1 U729 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n1223), .Y(n572) );
  MUX2X1 U730 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n1222), .Y(n571) );
  MUX2X1 U731 ( .B(n570), .A(n567), .S(n1189), .Y(n581) );
  MUX2X1 U732 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n1223), .Y(n575) );
  MUX2X1 U733 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n1222), .Y(n574) );
  MUX2X1 U734 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n1211), .Y(n578) );
  MUX2X1 U735 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n1213), .Y(n577) );
  MUX2X1 U736 ( .B(n576), .A(n573), .S(n1189), .Y(n580) );
  MUX2X1 U737 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n1223), .Y(n584) );
  MUX2X1 U738 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n1218), .Y(n583) );
  MUX2X1 U739 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n1222), .Y(n587) );
  MUX2X1 U740 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n1222), .Y(n586) );
  MUX2X1 U741 ( .B(n585), .A(n582), .S(n1189), .Y(n596) );
  MUX2X1 U742 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n1223), .Y(n590) );
  MUX2X1 U743 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n1223), .Y(n589) );
  MUX2X1 U744 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n1223), .Y(n593) );
  MUX2X1 U745 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n1223), .Y(n592) );
  MUX2X1 U746 ( .B(n591), .A(n588), .S(n1189), .Y(n595) );
  MUX2X1 U747 ( .B(n594), .A(n579), .S(n1185), .Y(n1182) );
  MUX2X1 U748 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n1223), .Y(n599) );
  MUX2X1 U749 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n1223), .Y(n598) );
  MUX2X1 U750 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n1223), .Y(n602) );
  MUX2X1 U751 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n1223), .Y(n601) );
  MUX2X1 U752 ( .B(n600), .A(n597), .S(n1189), .Y(n611) );
  MUX2X1 U753 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n1223), .Y(n605) );
  MUX2X1 U754 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n1223), .Y(n604) );
  MUX2X1 U755 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n1223), .Y(n608) );
  MUX2X1 U756 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n1223), .Y(n607) );
  MUX2X1 U757 ( .B(n606), .A(n603), .S(n1189), .Y(n610) );
  MUX2X1 U758 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n1223), .Y(n614) );
  MUX2X1 U759 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n1222), .Y(n613) );
  MUX2X1 U760 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n1218), .Y(n617) );
  MUX2X1 U761 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n1222), .Y(n616) );
  MUX2X1 U762 ( .B(n615), .A(n612), .S(n1189), .Y(n626) );
  MUX2X1 U763 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n1218), .Y(n620) );
  MUX2X1 U764 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n1223), .Y(n619) );
  MUX2X1 U765 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n1213), .Y(n623) );
  MUX2X1 U766 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n1218), .Y(n622) );
  MUX2X1 U767 ( .B(n621), .A(n618), .S(n1189), .Y(n625) );
  MUX2X1 U768 ( .B(n624), .A(n609), .S(n1185), .Y(n1183) );
  MUX2X1 U769 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n1211), .Y(n629) );
  MUX2X1 U770 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n1218), .Y(n628) );
  MUX2X1 U771 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n1211), .Y(n632) );
  MUX2X1 U772 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n1213), .Y(n631) );
  MUX2X1 U773 ( .B(n630), .A(n627), .S(n1192), .Y(n641) );
  MUX2X1 U774 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n1216), .Y(n635) );
  MUX2X1 U775 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n1218), .Y(n634) );
  MUX2X1 U776 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n1222), .Y(n638) );
  MUX2X1 U777 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n1221), .Y(n637) );
  MUX2X1 U778 ( .B(n636), .A(n633), .S(n1190), .Y(n640) );
  MUX2X1 U779 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n1218), .Y(n644) );
  MUX2X1 U780 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n1218), .Y(n643) );
  MUX2X1 U781 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n1223), .Y(n647) );
  MUX2X1 U782 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n1219), .Y(n646) );
  MUX2X1 U783 ( .B(n645), .A(n642), .S(n1190), .Y(n1168) );
  MUX2X1 U784 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n1223), .Y(n650) );
  MUX2X1 U785 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n1213), .Y(n649) );
  MUX2X1 U786 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n1218), .Y(n1165) );
  MUX2X1 U787 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n1216), .Y(n1164) );
  MUX2X1 U788 ( .B(n1163), .A(n648), .S(n1189), .Y(n1167) );
  MUX2X1 U789 ( .B(n1166), .A(n639), .S(n1185), .Y(n1184) );
  INVX1 U790 ( .A(N12), .Y(n1312) );
  INVX1 U791 ( .A(N11), .Y(n1310) );
  INVX1 U792 ( .A(write), .Y(n1226) );
  INVX1 U793 ( .A(n1226), .Y(n1227) );
  INVX1 U794 ( .A(N10), .Y(n1308) );
  INVX8 U795 ( .A(n1273), .Y(n1271) );
  INVX8 U796 ( .A(n62), .Y(n1275) );
  INVX8 U797 ( .A(n62), .Y(n1276) );
  INVX8 U798 ( .A(n65), .Y(n1277) );
  INVX8 U799 ( .A(n65), .Y(n1278) );
  INVX8 U800 ( .A(n66), .Y(n1279) );
  INVX8 U801 ( .A(n66), .Y(n1280) );
  INVX8 U802 ( .A(n67), .Y(n1281) );
  INVX8 U803 ( .A(n67), .Y(n1282) );
  INVX8 U804 ( .A(n68), .Y(n1283) );
  INVX8 U805 ( .A(n68), .Y(n1284) );
  INVX8 U806 ( .A(n69), .Y(n1285) );
  INVX8 U807 ( .A(n69), .Y(n1286) );
  INVX8 U808 ( .A(n70), .Y(n1287) );
  INVX8 U809 ( .A(n70), .Y(n1288) );
  INVX8 U810 ( .A(n71), .Y(n1289) );
  INVX8 U811 ( .A(n71), .Y(n1290) );
  INVX8 U812 ( .A(n72), .Y(n1291) );
  INVX8 U813 ( .A(n72), .Y(n1292) );
  INVX8 U814 ( .A(n73), .Y(n1293) );
  INVX8 U815 ( .A(n73), .Y(n1294) );
  INVX8 U816 ( .A(n74), .Y(n1295) );
  INVX8 U817 ( .A(n74), .Y(n1296) );
  INVX8 U818 ( .A(n75), .Y(n1297) );
  INVX8 U819 ( .A(n75), .Y(n1298) );
  INVX8 U820 ( .A(n76), .Y(n1299) );
  INVX8 U821 ( .A(n76), .Y(n1300) );
  INVX8 U822 ( .A(n77), .Y(n1301) );
  INVX8 U823 ( .A(n77), .Y(n1302) );
  INVX8 U824 ( .A(n78), .Y(n1303) );
  INVX8 U825 ( .A(n78), .Y(n1304) );
  INVX8 U826 ( .A(n79), .Y(n1305) );
  INVX8 U827 ( .A(n79), .Y(n1306) );
  OR2X2 U828 ( .A(write), .B(rst), .Y(n1316) );
  AND2X2 U829 ( .A(n20), .B(N32), .Y(\data_out<0> ) );
  AND2X2 U830 ( .A(n20), .B(N31), .Y(\data_out<1> ) );
  AND2X2 U831 ( .A(n1317), .B(N30), .Y(\data_out<2> ) );
  AND2X2 U832 ( .A(n20), .B(N29), .Y(\data_out<3> ) );
  AND2X2 U833 ( .A(n21), .B(N28), .Y(\data_out<4> ) );
  AND2X2 U834 ( .A(n20), .B(N27), .Y(\data_out<5> ) );
  AND2X2 U835 ( .A(N26), .B(n1317), .Y(\data_out<6> ) );
  AND2X2 U836 ( .A(n21), .B(N25), .Y(\data_out<7> ) );
  AND2X2 U837 ( .A(n20), .B(N24), .Y(\data_out<8> ) );
  AND2X2 U838 ( .A(n21), .B(N23), .Y(\data_out<9> ) );
  AND2X2 U839 ( .A(n21), .B(N22), .Y(\data_out<10> ) );
  AND2X2 U840 ( .A(n21), .B(N21), .Y(\data_out<11> ) );
  AND2X2 U841 ( .A(n21), .B(N20), .Y(\data_out<12> ) );
  AND2X2 U842 ( .A(n20), .B(N19), .Y(\data_out<13> ) );
  AND2X2 U843 ( .A(n21), .B(N18), .Y(\data_out<14> ) );
  AND2X2 U844 ( .A(n20), .B(N17), .Y(\data_out<15> ) );
  NAND2X1 U845 ( .A(\mem<31><0> ), .B(n1228), .Y(n1318) );
  OAI21X1 U846 ( .A(n121), .B(n1275), .C(n1318), .Y(n651) );
  NAND2X1 U847 ( .A(\mem<31><1> ), .B(n1229), .Y(n1319) );
  OAI21X1 U848 ( .A(n1278), .B(n121), .C(n1319), .Y(n652) );
  NAND2X1 U849 ( .A(\mem<31><2> ), .B(n1228), .Y(n1320) );
  OAI21X1 U850 ( .A(n1280), .B(n121), .C(n1320), .Y(n653) );
  NAND2X1 U851 ( .A(\mem<31><3> ), .B(n11), .Y(n1321) );
  OAI21X1 U852 ( .A(n1282), .B(n121), .C(n1321), .Y(n654) );
  NAND2X1 U853 ( .A(\mem<31><4> ), .B(n1229), .Y(n1322) );
  OAI21X1 U854 ( .A(n1284), .B(n121), .C(n1322), .Y(n655) );
  NAND2X1 U855 ( .A(\mem<31><5> ), .B(n1228), .Y(n1323) );
  OAI21X1 U856 ( .A(n1286), .B(n121), .C(n1323), .Y(n656) );
  NAND2X1 U857 ( .A(\mem<31><6> ), .B(n11), .Y(n1324) );
  OAI21X1 U858 ( .A(n1288), .B(n121), .C(n1324), .Y(n657) );
  NAND2X1 U859 ( .A(\mem<31><7> ), .B(n1229), .Y(n1325) );
  OAI21X1 U860 ( .A(n1290), .B(n121), .C(n1325), .Y(n658) );
  NAND2X1 U861 ( .A(\mem<31><8> ), .B(n1228), .Y(n1326) );
  OAI21X1 U862 ( .A(n1292), .B(n121), .C(n1326), .Y(n659) );
  NAND2X1 U863 ( .A(\mem<31><9> ), .B(n11), .Y(n1327) );
  OAI21X1 U864 ( .A(n1294), .B(n121), .C(n1327), .Y(n660) );
  NAND2X1 U865 ( .A(\mem<31><10> ), .B(n1229), .Y(n1328) );
  OAI21X1 U866 ( .A(n1296), .B(n121), .C(n1328), .Y(n661) );
  NAND2X1 U867 ( .A(\mem<31><11> ), .B(n1228), .Y(n1329) );
  OAI21X1 U868 ( .A(n1298), .B(n121), .C(n1329), .Y(n662) );
  NAND2X1 U869 ( .A(\mem<31><12> ), .B(n11), .Y(n1330) );
  OAI21X1 U870 ( .A(n1300), .B(n121), .C(n1330), .Y(n663) );
  NAND2X1 U871 ( .A(\mem<31><13> ), .B(n1229), .Y(n1331) );
  OAI21X1 U872 ( .A(n1302), .B(n121), .C(n1331), .Y(n664) );
  NAND2X1 U873 ( .A(\mem<31><14> ), .B(n1228), .Y(n1332) );
  OAI21X1 U874 ( .A(n1304), .B(n121), .C(n1332), .Y(n665) );
  NAND2X1 U875 ( .A(\mem<31><15> ), .B(n11), .Y(n1333) );
  OAI21X1 U876 ( .A(n1306), .B(n121), .C(n1333), .Y(n666) );
  NAND2X1 U877 ( .A(\mem<30><0> ), .B(n1230), .Y(n1334) );
  OAI21X1 U878 ( .A(n123), .B(n1275), .C(n1334), .Y(n667) );
  NAND2X1 U879 ( .A(\mem<30><1> ), .B(n10), .Y(n1335) );
  OAI21X1 U880 ( .A(n123), .B(n1278), .C(n1335), .Y(n668) );
  NAND2X1 U881 ( .A(\mem<30><2> ), .B(n1231), .Y(n1336) );
  OAI21X1 U882 ( .A(n123), .B(n1280), .C(n1336), .Y(n669) );
  NAND2X1 U883 ( .A(\mem<30><3> ), .B(n1230), .Y(n1337) );
  OAI21X1 U884 ( .A(n123), .B(n1282), .C(n1337), .Y(n670) );
  NAND2X1 U885 ( .A(\mem<30><4> ), .B(n10), .Y(n1338) );
  OAI21X1 U886 ( .A(n123), .B(n1284), .C(n1338), .Y(n671) );
  NAND2X1 U887 ( .A(\mem<30><5> ), .B(n1231), .Y(n1339) );
  OAI21X1 U888 ( .A(n123), .B(n1286), .C(n1339), .Y(n672) );
  NAND2X1 U889 ( .A(\mem<30><6> ), .B(n1230), .Y(n1340) );
  OAI21X1 U890 ( .A(n123), .B(n1288), .C(n1340), .Y(n673) );
  NAND2X1 U891 ( .A(\mem<30><7> ), .B(n10), .Y(n1341) );
  OAI21X1 U892 ( .A(n123), .B(n1290), .C(n1341), .Y(n674) );
  NAND2X1 U893 ( .A(\mem<30><8> ), .B(n1231), .Y(n1342) );
  OAI21X1 U894 ( .A(n123), .B(n1291), .C(n1342), .Y(n675) );
  NAND2X1 U895 ( .A(\mem<30><9> ), .B(n1230), .Y(n1343) );
  OAI21X1 U896 ( .A(n123), .B(n1293), .C(n1343), .Y(n676) );
  NAND2X1 U897 ( .A(\mem<30><10> ), .B(n10), .Y(n1344) );
  OAI21X1 U898 ( .A(n123), .B(n1295), .C(n1344), .Y(n677) );
  NAND2X1 U899 ( .A(\mem<30><11> ), .B(n1231), .Y(n1345) );
  OAI21X1 U900 ( .A(n123), .B(n1297), .C(n1345), .Y(n678) );
  NAND2X1 U901 ( .A(\mem<30><12> ), .B(n1230), .Y(n1346) );
  OAI21X1 U902 ( .A(n123), .B(n1299), .C(n1346), .Y(n679) );
  NAND2X1 U903 ( .A(\mem<30><13> ), .B(n10), .Y(n1347) );
  OAI21X1 U904 ( .A(n123), .B(n1301), .C(n1347), .Y(n680) );
  NAND2X1 U905 ( .A(\mem<30><14> ), .B(n1231), .Y(n1348) );
  OAI21X1 U906 ( .A(n123), .B(n1303), .C(n1348), .Y(n681) );
  NAND2X1 U907 ( .A(\mem<30><15> ), .B(n1230), .Y(n1349) );
  OAI21X1 U908 ( .A(n123), .B(n1305), .C(n1349), .Y(n682) );
  NAND3X1 U909 ( .A(n1219), .B(n1311), .C(n1310), .Y(n1350) );
  NAND2X1 U910 ( .A(\mem<29><0> ), .B(n1232), .Y(n1351) );
  OAI21X1 U911 ( .A(n125), .B(n1275), .C(n1351), .Y(n683) );
  NAND2X1 U912 ( .A(\mem<29><1> ), .B(n9), .Y(n1352) );
  OAI21X1 U913 ( .A(n125), .B(n1277), .C(n1352), .Y(n684) );
  NAND2X1 U914 ( .A(\mem<29><2> ), .B(n1233), .Y(n1353) );
  OAI21X1 U915 ( .A(n125), .B(n1279), .C(n1353), .Y(n685) );
  NAND2X1 U916 ( .A(\mem<29><3> ), .B(n1232), .Y(n1354) );
  OAI21X1 U917 ( .A(n125), .B(n1281), .C(n1354), .Y(n686) );
  NAND2X1 U918 ( .A(\mem<29><4> ), .B(n9), .Y(n1355) );
  OAI21X1 U919 ( .A(n125), .B(n1283), .C(n1355), .Y(n687) );
  NAND2X1 U920 ( .A(\mem<29><5> ), .B(n1233), .Y(n1356) );
  OAI21X1 U921 ( .A(n125), .B(n1285), .C(n1356), .Y(n688) );
  NAND2X1 U922 ( .A(\mem<29><6> ), .B(n1232), .Y(n1357) );
  OAI21X1 U923 ( .A(n125), .B(n1287), .C(n1357), .Y(n689) );
  NAND2X1 U924 ( .A(\mem<29><7> ), .B(n9), .Y(n1358) );
  OAI21X1 U925 ( .A(n125), .B(n1289), .C(n1358), .Y(n690) );
  NAND2X1 U926 ( .A(\mem<29><8> ), .B(n1233), .Y(n1359) );
  OAI21X1 U927 ( .A(n125), .B(n1292), .C(n1359), .Y(n691) );
  NAND2X1 U928 ( .A(\mem<29><9> ), .B(n1232), .Y(n1360) );
  OAI21X1 U929 ( .A(n125), .B(n1294), .C(n1360), .Y(n692) );
  NAND2X1 U930 ( .A(\mem<29><10> ), .B(n9), .Y(n1361) );
  OAI21X1 U931 ( .A(n125), .B(n1296), .C(n1361), .Y(n693) );
  NAND2X1 U932 ( .A(\mem<29><11> ), .B(n1233), .Y(n1362) );
  OAI21X1 U933 ( .A(n125), .B(n1298), .C(n1362), .Y(n694) );
  NAND2X1 U934 ( .A(\mem<29><12> ), .B(n1232), .Y(n1363) );
  OAI21X1 U935 ( .A(n125), .B(n1300), .C(n1363), .Y(n695) );
  NAND2X1 U936 ( .A(\mem<29><13> ), .B(n9), .Y(n1364) );
  OAI21X1 U937 ( .A(n125), .B(n1302), .C(n1364), .Y(n696) );
  NAND2X1 U938 ( .A(\mem<29><14> ), .B(n1233), .Y(n1365) );
  OAI21X1 U939 ( .A(n125), .B(n1304), .C(n1365), .Y(n697) );
  NAND2X1 U940 ( .A(\mem<29><15> ), .B(n1232), .Y(n1366) );
  OAI21X1 U941 ( .A(n125), .B(n1306), .C(n1366), .Y(n698) );
  NAND3X1 U942 ( .A(n1311), .B(n1310), .C(n1308), .Y(n1367) );
  NAND2X1 U943 ( .A(\mem<28><0> ), .B(n1234), .Y(n1368) );
  OAI21X1 U944 ( .A(n127), .B(n1275), .C(n1368), .Y(n699) );
  NAND2X1 U945 ( .A(\mem<28><1> ), .B(n8), .Y(n1369) );
  OAI21X1 U946 ( .A(n127), .B(n1278), .C(n1369), .Y(n700) );
  NAND2X1 U947 ( .A(\mem<28><2> ), .B(n1235), .Y(n1370) );
  OAI21X1 U948 ( .A(n127), .B(n1280), .C(n1370), .Y(n701) );
  NAND2X1 U949 ( .A(\mem<28><3> ), .B(n1234), .Y(n1371) );
  OAI21X1 U950 ( .A(n127), .B(n1282), .C(n1371), .Y(n702) );
  NAND2X1 U951 ( .A(\mem<28><4> ), .B(n8), .Y(n1372) );
  OAI21X1 U952 ( .A(n127), .B(n1284), .C(n1372), .Y(n703) );
  NAND2X1 U953 ( .A(\mem<28><5> ), .B(n1235), .Y(n1373) );
  OAI21X1 U954 ( .A(n127), .B(n1286), .C(n1373), .Y(n704) );
  NAND2X1 U955 ( .A(\mem<28><6> ), .B(n1234), .Y(n1374) );
  OAI21X1 U956 ( .A(n127), .B(n1288), .C(n1374), .Y(n705) );
  NAND2X1 U957 ( .A(\mem<28><7> ), .B(n8), .Y(n1375) );
  OAI21X1 U958 ( .A(n127), .B(n1290), .C(n1375), .Y(n706) );
  NAND2X1 U959 ( .A(\mem<28><8> ), .B(n1235), .Y(n1376) );
  OAI21X1 U960 ( .A(n127), .B(n1291), .C(n1376), .Y(n707) );
  NAND2X1 U961 ( .A(\mem<28><9> ), .B(n1234), .Y(n1377) );
  OAI21X1 U962 ( .A(n127), .B(n1293), .C(n1377), .Y(n708) );
  NAND2X1 U963 ( .A(\mem<28><10> ), .B(n8), .Y(n1378) );
  OAI21X1 U964 ( .A(n127), .B(n1295), .C(n1378), .Y(n709) );
  NAND2X1 U965 ( .A(\mem<28><11> ), .B(n1235), .Y(n1379) );
  OAI21X1 U966 ( .A(n127), .B(n1297), .C(n1379), .Y(n710) );
  NAND2X1 U967 ( .A(\mem<28><12> ), .B(n1234), .Y(n1380) );
  OAI21X1 U968 ( .A(n127), .B(n1299), .C(n1380), .Y(n711) );
  NAND2X1 U969 ( .A(\mem<28><13> ), .B(n8), .Y(n1381) );
  OAI21X1 U970 ( .A(n127), .B(n1301), .C(n1381), .Y(n712) );
  NAND2X1 U971 ( .A(\mem<28><14> ), .B(n1235), .Y(n1382) );
  OAI21X1 U972 ( .A(n127), .B(n1303), .C(n1382), .Y(n713) );
  NAND2X1 U973 ( .A(\mem<28><15> ), .B(n1234), .Y(n1383) );
  OAI21X1 U974 ( .A(n127), .B(n1305), .C(n1383), .Y(n714) );
  NAND3X1 U975 ( .A(n1212), .B(n1309), .C(n1312), .Y(n1384) );
  NAND2X1 U976 ( .A(\mem<27><0> ), .B(n1236), .Y(n1385) );
  OAI21X1 U977 ( .A(n129), .B(n1275), .C(n1385), .Y(n715) );
  NAND2X1 U978 ( .A(\mem<27><1> ), .B(n7), .Y(n1386) );
  OAI21X1 U979 ( .A(n129), .B(n1277), .C(n1386), .Y(n716) );
  NAND2X1 U980 ( .A(\mem<27><2> ), .B(n1237), .Y(n1387) );
  OAI21X1 U981 ( .A(n129), .B(n1279), .C(n1387), .Y(n717) );
  NAND2X1 U982 ( .A(\mem<27><3> ), .B(n1236), .Y(n1388) );
  OAI21X1 U983 ( .A(n129), .B(n1281), .C(n1388), .Y(n718) );
  NAND2X1 U984 ( .A(\mem<27><4> ), .B(n7), .Y(n1389) );
  OAI21X1 U985 ( .A(n129), .B(n1283), .C(n1389), .Y(n719) );
  NAND2X1 U986 ( .A(\mem<27><5> ), .B(n1237), .Y(n1390) );
  OAI21X1 U987 ( .A(n129), .B(n1285), .C(n1390), .Y(n720) );
  NAND2X1 U988 ( .A(\mem<27><6> ), .B(n1236), .Y(n1391) );
  OAI21X1 U989 ( .A(n129), .B(n1287), .C(n1391), .Y(n721) );
  NAND2X1 U990 ( .A(\mem<27><7> ), .B(n7), .Y(n1392) );
  OAI21X1 U991 ( .A(n129), .B(n1289), .C(n1392), .Y(n722) );
  NAND2X1 U992 ( .A(\mem<27><8> ), .B(n1237), .Y(n1393) );
  OAI21X1 U993 ( .A(n129), .B(n1292), .C(n1393), .Y(n723) );
  NAND2X1 U994 ( .A(\mem<27><9> ), .B(n1236), .Y(n1394) );
  OAI21X1 U995 ( .A(n129), .B(n1294), .C(n1394), .Y(n724) );
  NAND2X1 U996 ( .A(\mem<27><10> ), .B(n7), .Y(n1395) );
  OAI21X1 U997 ( .A(n129), .B(n1296), .C(n1395), .Y(n725) );
  NAND2X1 U998 ( .A(\mem<27><11> ), .B(n1237), .Y(n1396) );
  OAI21X1 U999 ( .A(n129), .B(n1298), .C(n1396), .Y(n726) );
  NAND2X1 U1000 ( .A(\mem<27><12> ), .B(n1236), .Y(n1397) );
  OAI21X1 U1001 ( .A(n129), .B(n1300), .C(n1397), .Y(n727) );
  NAND2X1 U1002 ( .A(\mem<27><13> ), .B(n7), .Y(n1398) );
  OAI21X1 U1003 ( .A(n129), .B(n1302), .C(n1398), .Y(n728) );
  NAND2X1 U1004 ( .A(\mem<27><14> ), .B(n1237), .Y(n1399) );
  OAI21X1 U1005 ( .A(n129), .B(n1304), .C(n1399), .Y(n729) );
  NAND2X1 U1006 ( .A(\mem<27><15> ), .B(n1236), .Y(n1400) );
  OAI21X1 U1007 ( .A(n129), .B(n1306), .C(n1400), .Y(n730) );
  NAND3X1 U1008 ( .A(n1312), .B(n1309), .C(n1308), .Y(n1401) );
  NAND2X1 U1009 ( .A(\mem<26><0> ), .B(n1238), .Y(n1402) );
  OAI21X1 U1010 ( .A(n131), .B(n1275), .C(n1402), .Y(n731) );
  NAND2X1 U1011 ( .A(\mem<26><1> ), .B(n6), .Y(n1403) );
  OAI21X1 U1012 ( .A(n131), .B(n1278), .C(n1403), .Y(n732) );
  NAND2X1 U1013 ( .A(\mem<26><2> ), .B(n1239), .Y(n1404) );
  OAI21X1 U1014 ( .A(n131), .B(n1280), .C(n1404), .Y(n733) );
  NAND2X1 U1015 ( .A(\mem<26><3> ), .B(n1238), .Y(n1405) );
  OAI21X1 U1016 ( .A(n131), .B(n1282), .C(n1405), .Y(n734) );
  NAND2X1 U1017 ( .A(\mem<26><4> ), .B(n6), .Y(n1406) );
  OAI21X1 U1018 ( .A(n131), .B(n1284), .C(n1406), .Y(n735) );
  NAND2X1 U1019 ( .A(\mem<26><5> ), .B(n1239), .Y(n1407) );
  OAI21X1 U1020 ( .A(n131), .B(n1286), .C(n1407), .Y(n736) );
  NAND2X1 U1021 ( .A(\mem<26><6> ), .B(n1238), .Y(n1408) );
  OAI21X1 U1022 ( .A(n131), .B(n1288), .C(n1408), .Y(n737) );
  NAND2X1 U1023 ( .A(\mem<26><7> ), .B(n6), .Y(n1409) );
  OAI21X1 U1024 ( .A(n131), .B(n1290), .C(n1409), .Y(n738) );
  NAND2X1 U1025 ( .A(\mem<26><8> ), .B(n1239), .Y(n1410) );
  OAI21X1 U1026 ( .A(n131), .B(n1291), .C(n1410), .Y(n739) );
  NAND2X1 U1027 ( .A(\mem<26><9> ), .B(n1238), .Y(n1411) );
  OAI21X1 U1028 ( .A(n131), .B(n1293), .C(n1411), .Y(n740) );
  NAND2X1 U1029 ( .A(\mem<26><10> ), .B(n6), .Y(n1412) );
  OAI21X1 U1030 ( .A(n131), .B(n1295), .C(n1412), .Y(n741) );
  NAND2X1 U1031 ( .A(\mem<26><11> ), .B(n1239), .Y(n1413) );
  OAI21X1 U1032 ( .A(n131), .B(n1297), .C(n1413), .Y(n742) );
  NAND2X1 U1033 ( .A(\mem<26><12> ), .B(n1238), .Y(n1414) );
  OAI21X1 U1034 ( .A(n131), .B(n1299), .C(n1414), .Y(n743) );
  NAND2X1 U1035 ( .A(\mem<26><13> ), .B(n6), .Y(n1415) );
  OAI21X1 U1036 ( .A(n131), .B(n1301), .C(n1415), .Y(n744) );
  NAND2X1 U1037 ( .A(\mem<26><14> ), .B(n1239), .Y(n1416) );
  OAI21X1 U1038 ( .A(n131), .B(n1303), .C(n1416), .Y(n745) );
  NAND2X1 U1039 ( .A(\mem<26><15> ), .B(n1238), .Y(n1417) );
  OAI21X1 U1040 ( .A(n131), .B(n1305), .C(n1417), .Y(n746) );
  NAND3X1 U1041 ( .A(n1210), .B(n1312), .C(n1310), .Y(n1418) );
  NAND2X1 U1042 ( .A(\mem<25><0> ), .B(n1240), .Y(n1419) );
  OAI21X1 U1043 ( .A(n133), .B(n1275), .C(n1419), .Y(n747) );
  NAND2X1 U1044 ( .A(\mem<25><1> ), .B(n5), .Y(n1420) );
  OAI21X1 U1045 ( .A(n133), .B(n1277), .C(n1420), .Y(n748) );
  NAND2X1 U1046 ( .A(\mem<25><2> ), .B(n1241), .Y(n1421) );
  OAI21X1 U1047 ( .A(n133), .B(n1279), .C(n1421), .Y(n749) );
  NAND2X1 U1048 ( .A(\mem<25><3> ), .B(n1240), .Y(n1422) );
  OAI21X1 U1049 ( .A(n133), .B(n1281), .C(n1422), .Y(n750) );
  NAND2X1 U1050 ( .A(\mem<25><4> ), .B(n5), .Y(n1423) );
  OAI21X1 U1051 ( .A(n133), .B(n1283), .C(n1423), .Y(n751) );
  NAND2X1 U1052 ( .A(\mem<25><5> ), .B(n1241), .Y(n1424) );
  OAI21X1 U1053 ( .A(n133), .B(n1285), .C(n1424), .Y(n752) );
  NAND2X1 U1054 ( .A(\mem<25><6> ), .B(n1240), .Y(n1425) );
  OAI21X1 U1055 ( .A(n133), .B(n1287), .C(n1425), .Y(n753) );
  NAND2X1 U1056 ( .A(\mem<25><7> ), .B(n5), .Y(n1426) );
  OAI21X1 U1057 ( .A(n133), .B(n1289), .C(n1426), .Y(n754) );
  NAND2X1 U1058 ( .A(\mem<25><8> ), .B(n1241), .Y(n1427) );
  OAI21X1 U1059 ( .A(n133), .B(n1292), .C(n1427), .Y(n755) );
  NAND2X1 U1060 ( .A(\mem<25><9> ), .B(n1240), .Y(n1428) );
  OAI21X1 U1061 ( .A(n133), .B(n1294), .C(n1428), .Y(n756) );
  NAND2X1 U1062 ( .A(\mem<25><10> ), .B(n5), .Y(n1429) );
  OAI21X1 U1063 ( .A(n133), .B(n1296), .C(n1429), .Y(n757) );
  NAND2X1 U1064 ( .A(\mem<25><11> ), .B(n1241), .Y(n1430) );
  OAI21X1 U1065 ( .A(n133), .B(n1298), .C(n1430), .Y(n758) );
  NAND2X1 U1066 ( .A(\mem<25><12> ), .B(n1240), .Y(n1431) );
  OAI21X1 U1067 ( .A(n133), .B(n1300), .C(n1431), .Y(n759) );
  NAND2X1 U1068 ( .A(\mem<25><13> ), .B(n5), .Y(n1432) );
  OAI21X1 U1069 ( .A(n133), .B(n1302), .C(n1432), .Y(n760) );
  NAND2X1 U1070 ( .A(\mem<25><14> ), .B(n1241), .Y(n1433) );
  OAI21X1 U1071 ( .A(n133), .B(n1304), .C(n1433), .Y(n761) );
  NAND2X1 U1072 ( .A(\mem<25><15> ), .B(n1240), .Y(n1434) );
  OAI21X1 U1073 ( .A(n133), .B(n1306), .C(n1434), .Y(n762) );
  NOR3X1 U1074 ( .A(n1210), .B(n1309), .C(n1311), .Y(n1828) );
  NAND2X1 U1075 ( .A(\mem<24><0> ), .B(n1243), .Y(n1435) );
  OAI21X1 U1076 ( .A(n1242), .B(n1275), .C(n1435), .Y(n763) );
  NAND2X1 U1077 ( .A(\mem<24><1> ), .B(n12), .Y(n1436) );
  OAI21X1 U1078 ( .A(n1242), .B(n1277), .C(n1436), .Y(n764) );
  NAND2X1 U1079 ( .A(\mem<24><2> ), .B(n1244), .Y(n1437) );
  OAI21X1 U1080 ( .A(n1242), .B(n1279), .C(n1437), .Y(n765) );
  NAND2X1 U1081 ( .A(\mem<24><3> ), .B(n1243), .Y(n1438) );
  OAI21X1 U1082 ( .A(n1242), .B(n1281), .C(n1438), .Y(n766) );
  NAND2X1 U1083 ( .A(\mem<24><4> ), .B(n12), .Y(n1439) );
  OAI21X1 U1084 ( .A(n1242), .B(n1283), .C(n1439), .Y(n767) );
  NAND2X1 U1085 ( .A(\mem<24><5> ), .B(n1244), .Y(n1440) );
  OAI21X1 U1086 ( .A(n1242), .B(n1285), .C(n1440), .Y(n768) );
  NAND2X1 U1087 ( .A(\mem<24><6> ), .B(n1243), .Y(n1441) );
  OAI21X1 U1088 ( .A(n1242), .B(n1287), .C(n1441), .Y(n769) );
  NAND2X1 U1089 ( .A(\mem<24><7> ), .B(n12), .Y(n1442) );
  OAI21X1 U1090 ( .A(n1242), .B(n1289), .C(n1442), .Y(n770) );
  NAND2X1 U1091 ( .A(\mem<24><8> ), .B(n1244), .Y(n1443) );
  OAI21X1 U1092 ( .A(n1242), .B(n1291), .C(n1443), .Y(n771) );
  NAND2X1 U1093 ( .A(\mem<24><9> ), .B(n1243), .Y(n1444) );
  OAI21X1 U1094 ( .A(n1242), .B(n1293), .C(n1444), .Y(n772) );
  NAND2X1 U1095 ( .A(\mem<24><10> ), .B(n1243), .Y(n1445) );
  OAI21X1 U1096 ( .A(n1242), .B(n1295), .C(n1445), .Y(n773) );
  NAND2X1 U1097 ( .A(\mem<24><11> ), .B(n12), .Y(n1446) );
  OAI21X1 U1098 ( .A(n1242), .B(n1297), .C(n1446), .Y(n774) );
  NAND2X1 U1099 ( .A(\mem<24><12> ), .B(n12), .Y(n1447) );
  OAI21X1 U1100 ( .A(n1242), .B(n1299), .C(n1447), .Y(n775) );
  NAND2X1 U1101 ( .A(\mem<24><13> ), .B(n1244), .Y(n1448) );
  OAI21X1 U1102 ( .A(n1242), .B(n1301), .C(n1448), .Y(n776) );
  NAND2X1 U1103 ( .A(\mem<24><14> ), .B(n1244), .Y(n1449) );
  OAI21X1 U1104 ( .A(n1242), .B(n1303), .C(n1449), .Y(n777) );
  NAND2X1 U1105 ( .A(\mem<24><15> ), .B(n1243), .Y(n1450) );
  OAI21X1 U1106 ( .A(n1242), .B(n1305), .C(n1450), .Y(n778) );
  NAND2X1 U1107 ( .A(\mem<23><0> ), .B(n1245), .Y(n1451) );
  OAI21X1 U1108 ( .A(n135), .B(n1275), .C(n1451), .Y(n779) );
  NAND2X1 U1109 ( .A(\mem<23><1> ), .B(n4), .Y(n1452) );
  OAI21X1 U1110 ( .A(n135), .B(n1278), .C(n1452), .Y(n780) );
  NAND2X1 U1111 ( .A(\mem<23><2> ), .B(n1246), .Y(n1453) );
  OAI21X1 U1112 ( .A(n135), .B(n1280), .C(n1453), .Y(n781) );
  NAND2X1 U1113 ( .A(\mem<23><3> ), .B(n1245), .Y(n1454) );
  OAI21X1 U1114 ( .A(n135), .B(n1282), .C(n1454), .Y(n782) );
  NAND2X1 U1115 ( .A(\mem<23><4> ), .B(n4), .Y(n1455) );
  OAI21X1 U1116 ( .A(n135), .B(n1284), .C(n1455), .Y(n783) );
  NAND2X1 U1117 ( .A(\mem<23><5> ), .B(n1246), .Y(n1456) );
  OAI21X1 U1118 ( .A(n135), .B(n1286), .C(n1456), .Y(n784) );
  NAND2X1 U1119 ( .A(\mem<23><6> ), .B(n1245), .Y(n1457) );
  OAI21X1 U1120 ( .A(n135), .B(n1288), .C(n1457), .Y(n785) );
  NAND2X1 U1121 ( .A(\mem<23><7> ), .B(n4), .Y(n1458) );
  OAI21X1 U1122 ( .A(n135), .B(n1290), .C(n1458), .Y(n786) );
  NAND2X1 U1123 ( .A(\mem<23><8> ), .B(n1246), .Y(n1459) );
  OAI21X1 U1124 ( .A(n135), .B(n1292), .C(n1459), .Y(n787) );
  NAND2X1 U1125 ( .A(\mem<23><9> ), .B(n1245), .Y(n1460) );
  OAI21X1 U1126 ( .A(n135), .B(n1294), .C(n1460), .Y(n788) );
  NAND2X1 U1127 ( .A(\mem<23><10> ), .B(n4), .Y(n1461) );
  OAI21X1 U1128 ( .A(n135), .B(n1296), .C(n1461), .Y(n789) );
  NAND2X1 U1129 ( .A(\mem<23><11> ), .B(n1246), .Y(n1462) );
  OAI21X1 U1130 ( .A(n135), .B(n1298), .C(n1462), .Y(n790) );
  NAND2X1 U1131 ( .A(\mem<23><12> ), .B(n1245), .Y(n1463) );
  OAI21X1 U1132 ( .A(n135), .B(n1300), .C(n1463), .Y(n791) );
  NAND2X1 U1133 ( .A(\mem<23><13> ), .B(n4), .Y(n1464) );
  OAI21X1 U1134 ( .A(n135), .B(n1302), .C(n1464), .Y(n792) );
  NAND2X1 U1135 ( .A(\mem<23><14> ), .B(n1246), .Y(n1465) );
  OAI21X1 U1136 ( .A(n135), .B(n1304), .C(n1465), .Y(n793) );
  NAND2X1 U1137 ( .A(\mem<23><15> ), .B(n1245), .Y(n1466) );
  OAI21X1 U1138 ( .A(n135), .B(n1306), .C(n1466), .Y(n794) );
  NAND2X1 U1139 ( .A(\mem<22><0> ), .B(n1247), .Y(n1467) );
  OAI21X1 U1140 ( .A(n137), .B(n1275), .C(n1467), .Y(n795) );
  NAND2X1 U1141 ( .A(\mem<22><1> ), .B(n3), .Y(n1468) );
  OAI21X1 U1142 ( .A(n137), .B(n1278), .C(n1468), .Y(n796) );
  NAND2X1 U1143 ( .A(\mem<22><2> ), .B(n1248), .Y(n1469) );
  OAI21X1 U1144 ( .A(n137), .B(n1280), .C(n1469), .Y(n797) );
  NAND2X1 U1145 ( .A(\mem<22><3> ), .B(n1247), .Y(n1470) );
  OAI21X1 U1146 ( .A(n137), .B(n1282), .C(n1470), .Y(n798) );
  NAND2X1 U1147 ( .A(\mem<22><4> ), .B(n3), .Y(n1471) );
  OAI21X1 U1148 ( .A(n137), .B(n1284), .C(n1471), .Y(n799) );
  NAND2X1 U1149 ( .A(\mem<22><5> ), .B(n1248), .Y(n1472) );
  OAI21X1 U1150 ( .A(n137), .B(n1286), .C(n1472), .Y(n800) );
  NAND2X1 U1151 ( .A(\mem<22><6> ), .B(n1247), .Y(n1473) );
  OAI21X1 U1152 ( .A(n137), .B(n1288), .C(n1473), .Y(n801) );
  NAND2X1 U1153 ( .A(\mem<22><7> ), .B(n3), .Y(n1474) );
  OAI21X1 U1154 ( .A(n137), .B(n1290), .C(n1474), .Y(n802) );
  NAND2X1 U1155 ( .A(\mem<22><8> ), .B(n1248), .Y(n1475) );
  OAI21X1 U1156 ( .A(n137), .B(n1292), .C(n1475), .Y(n803) );
  NAND2X1 U1157 ( .A(\mem<22><9> ), .B(n1247), .Y(n1476) );
  OAI21X1 U1158 ( .A(n137), .B(n1294), .C(n1476), .Y(n804) );
  NAND2X1 U1159 ( .A(\mem<22><10> ), .B(n3), .Y(n1477) );
  OAI21X1 U1160 ( .A(n137), .B(n1296), .C(n1477), .Y(n805) );
  NAND2X1 U1161 ( .A(\mem<22><11> ), .B(n1248), .Y(n1478) );
  OAI21X1 U1162 ( .A(n137), .B(n1298), .C(n1478), .Y(n806) );
  NAND2X1 U1163 ( .A(\mem<22><12> ), .B(n1247), .Y(n1479) );
  OAI21X1 U1164 ( .A(n137), .B(n1300), .C(n1479), .Y(n807) );
  NAND2X1 U1165 ( .A(\mem<22><13> ), .B(n3), .Y(n1480) );
  OAI21X1 U1166 ( .A(n137), .B(n1302), .C(n1480), .Y(n808) );
  NAND2X1 U1167 ( .A(\mem<22><14> ), .B(n1248), .Y(n1481) );
  OAI21X1 U1168 ( .A(n137), .B(n1304), .C(n1481), .Y(n809) );
  NAND2X1 U1169 ( .A(\mem<22><15> ), .B(n1247), .Y(n1482) );
  OAI21X1 U1170 ( .A(n137), .B(n1306), .C(n1482), .Y(n810) );
  NAND2X1 U1171 ( .A(\mem<21><0> ), .B(n1249), .Y(n1483) );
  OAI21X1 U1172 ( .A(n139), .B(n1275), .C(n1483), .Y(n811) );
  NAND2X1 U1173 ( .A(\mem<21><1> ), .B(n2), .Y(n1484) );
  OAI21X1 U1174 ( .A(n139), .B(n1278), .C(n1484), .Y(n812) );
  NAND2X1 U1175 ( .A(\mem<21><2> ), .B(n1250), .Y(n1485) );
  OAI21X1 U1177 ( .A(n139), .B(n1280), .C(n1485), .Y(n813) );
  NAND2X1 U1178 ( .A(\mem<21><3> ), .B(n1249), .Y(n1486) );
  OAI21X1 U1179 ( .A(n139), .B(n1282), .C(n1486), .Y(n814) );
  NAND2X1 U1180 ( .A(\mem<21><4> ), .B(n2), .Y(n1487) );
  OAI21X1 U1181 ( .A(n139), .B(n1284), .C(n1487), .Y(n815) );
  NAND2X1 U1182 ( .A(\mem<21><5> ), .B(n1250), .Y(n1488) );
  OAI21X1 U1183 ( .A(n139), .B(n1286), .C(n1488), .Y(n816) );
  NAND2X1 U1184 ( .A(\mem<21><6> ), .B(n1249), .Y(n1489) );
  OAI21X1 U1185 ( .A(n139), .B(n1288), .C(n1489), .Y(n817) );
  NAND2X1 U1186 ( .A(\mem<21><7> ), .B(n2), .Y(n1490) );
  OAI21X1 U1187 ( .A(n139), .B(n1290), .C(n1490), .Y(n818) );
  NAND2X1 U1188 ( .A(\mem<21><8> ), .B(n1250), .Y(n1491) );
  OAI21X1 U1189 ( .A(n139), .B(n1292), .C(n1491), .Y(n819) );
  NAND2X1 U1190 ( .A(\mem<21><9> ), .B(n1249), .Y(n1492) );
  OAI21X1 U1191 ( .A(n139), .B(n1294), .C(n1492), .Y(n820) );
  NAND2X1 U1192 ( .A(\mem<21><10> ), .B(n2), .Y(n1493) );
  OAI21X1 U1193 ( .A(n139), .B(n1296), .C(n1493), .Y(n821) );
  NAND2X1 U1194 ( .A(\mem<21><11> ), .B(n1250), .Y(n1494) );
  OAI21X1 U1195 ( .A(n139), .B(n1298), .C(n1494), .Y(n822) );
  NAND2X1 U1196 ( .A(\mem<21><12> ), .B(n1249), .Y(n1495) );
  OAI21X1 U1197 ( .A(n139), .B(n1300), .C(n1495), .Y(n823) );
  NAND2X1 U1198 ( .A(\mem<21><13> ), .B(n2), .Y(n1496) );
  OAI21X1 U1199 ( .A(n139), .B(n1302), .C(n1496), .Y(n824) );
  NAND2X1 U1200 ( .A(\mem<21><14> ), .B(n1250), .Y(n1497) );
  OAI21X1 U1201 ( .A(n139), .B(n1304), .C(n1497), .Y(n825) );
  NAND2X1 U1202 ( .A(\mem<21><15> ), .B(n1249), .Y(n1498) );
  OAI21X1 U1203 ( .A(n139), .B(n1306), .C(n1498), .Y(n826) );
  NAND2X1 U1204 ( .A(\mem<20><0> ), .B(n1252), .Y(n1499) );
  OAI21X1 U1205 ( .A(n141), .B(n1275), .C(n1499), .Y(n827) );
  NAND2X1 U1206 ( .A(\mem<20><1> ), .B(n1), .Y(n1500) );
  OAI21X1 U1207 ( .A(n141), .B(n1278), .C(n1500), .Y(n828) );
  NAND2X1 U1208 ( .A(\mem<20><2> ), .B(n1252), .Y(n1501) );
  OAI21X1 U1209 ( .A(n141), .B(n1280), .C(n1501), .Y(n829) );
  NAND2X1 U1210 ( .A(\mem<20><3> ), .B(n1), .Y(n1502) );
  OAI21X1 U1211 ( .A(n141), .B(n1282), .C(n1502), .Y(n830) );
  NAND2X1 U1212 ( .A(\mem<20><4> ), .B(n1252), .Y(n1503) );
  OAI21X1 U1213 ( .A(n141), .B(n1284), .C(n1503), .Y(n831) );
  NAND2X1 U1214 ( .A(\mem<20><5> ), .B(n1), .Y(n1504) );
  OAI21X1 U1215 ( .A(n141), .B(n1286), .C(n1504), .Y(n832) );
  NAND2X1 U1216 ( .A(\mem<20><6> ), .B(n1252), .Y(n1505) );
  OAI21X1 U1217 ( .A(n141), .B(n1288), .C(n1505), .Y(n833) );
  NAND2X1 U1218 ( .A(\mem<20><7> ), .B(n1), .Y(n1506) );
  OAI21X1 U1219 ( .A(n141), .B(n1290), .C(n1506), .Y(n834) );
  NAND2X1 U1220 ( .A(\mem<20><8> ), .B(n1252), .Y(n1507) );
  OAI21X1 U1221 ( .A(n141), .B(n1292), .C(n1507), .Y(n835) );
  NAND2X1 U1222 ( .A(\mem<20><9> ), .B(n1), .Y(n1508) );
  OAI21X1 U1223 ( .A(n141), .B(n1294), .C(n1508), .Y(n836) );
  NAND2X1 U1224 ( .A(\mem<20><10> ), .B(n1251), .Y(n1509) );
  OAI21X1 U1225 ( .A(n141), .B(n1296), .C(n1509), .Y(n837) );
  NAND2X1 U1226 ( .A(\mem<20><11> ), .B(n1251), .Y(n1510) );
  OAI21X1 U1227 ( .A(n141), .B(n1298), .C(n1510), .Y(n838) );
  NAND2X1 U1228 ( .A(\mem<20><12> ), .B(n1251), .Y(n1511) );
  OAI21X1 U1229 ( .A(n141), .B(n1300), .C(n1511), .Y(n839) );
  NAND2X1 U1230 ( .A(\mem<20><13> ), .B(n1251), .Y(n1512) );
  OAI21X1 U1231 ( .A(n141), .B(n1302), .C(n1512), .Y(n840) );
  NAND2X1 U1232 ( .A(\mem<20><14> ), .B(n1251), .Y(n1513) );
  OAI21X1 U1233 ( .A(n141), .B(n1304), .C(n1513), .Y(n841) );
  NAND2X1 U1234 ( .A(\mem<20><15> ), .B(n1251), .Y(n1514) );
  OAI21X1 U1235 ( .A(n141), .B(n1306), .C(n1514), .Y(n842) );
  NAND2X1 U1236 ( .A(\mem<19><0> ), .B(n23), .Y(n1515) );
  OAI21X1 U1237 ( .A(n143), .B(n1276), .C(n1515), .Y(n843) );
  NAND2X1 U1238 ( .A(\mem<19><1> ), .B(n23), .Y(n1516) );
  OAI21X1 U1239 ( .A(n143), .B(n1278), .C(n1516), .Y(n844) );
  NAND2X1 U1240 ( .A(\mem<19><2> ), .B(n23), .Y(n1517) );
  OAI21X1 U1241 ( .A(n143), .B(n1280), .C(n1517), .Y(n845) );
  NAND2X1 U1242 ( .A(\mem<19><3> ), .B(n23), .Y(n1518) );
  OAI21X1 U1243 ( .A(n143), .B(n1282), .C(n1518), .Y(n846) );
  NAND2X1 U1244 ( .A(\mem<19><4> ), .B(n23), .Y(n1519) );
  OAI21X1 U1245 ( .A(n143), .B(n1284), .C(n1519), .Y(n847) );
  NAND2X1 U1246 ( .A(\mem<19><5> ), .B(n23), .Y(n1520) );
  OAI21X1 U1247 ( .A(n143), .B(n1286), .C(n1520), .Y(n848) );
  NAND2X1 U1248 ( .A(\mem<19><6> ), .B(n23), .Y(n1521) );
  OAI21X1 U1249 ( .A(n143), .B(n1288), .C(n1521), .Y(n849) );
  NAND2X1 U1250 ( .A(\mem<19><7> ), .B(n23), .Y(n1522) );
  OAI21X1 U1251 ( .A(n143), .B(n1290), .C(n1522), .Y(n850) );
  NAND2X1 U1252 ( .A(\mem<19><8> ), .B(n23), .Y(n1523) );
  OAI21X1 U1253 ( .A(n143), .B(n1292), .C(n1523), .Y(n851) );
  NAND2X1 U1254 ( .A(\mem<19><9> ), .B(n23), .Y(n1524) );
  OAI21X1 U1255 ( .A(n143), .B(n1294), .C(n1524), .Y(n852) );
  NAND2X1 U1256 ( .A(\mem<19><10> ), .B(n23), .Y(n1525) );
  OAI21X1 U1257 ( .A(n143), .B(n1296), .C(n1525), .Y(n853) );
  NAND2X1 U1258 ( .A(\mem<19><11> ), .B(n23), .Y(n1526) );
  OAI21X1 U1259 ( .A(n143), .B(n1298), .C(n1526), .Y(n854) );
  NAND2X1 U1260 ( .A(\mem<19><12> ), .B(n23), .Y(n1527) );
  OAI21X1 U1261 ( .A(n143), .B(n1300), .C(n1527), .Y(n855) );
  NAND2X1 U1262 ( .A(\mem<19><13> ), .B(n23), .Y(n1528) );
  OAI21X1 U1263 ( .A(n143), .B(n1302), .C(n1528), .Y(n856) );
  NAND2X1 U1264 ( .A(\mem<19><14> ), .B(n23), .Y(n1529) );
  OAI21X1 U1265 ( .A(n143), .B(n1304), .C(n1529), .Y(n857) );
  NAND2X1 U1266 ( .A(\mem<19><15> ), .B(n23), .Y(n1530) );
  OAI21X1 U1267 ( .A(n143), .B(n1306), .C(n1530), .Y(n858) );
  NAND2X1 U1268 ( .A(\mem<18><0> ), .B(n25), .Y(n1531) );
  OAI21X1 U1269 ( .A(n145), .B(n1276), .C(n1531), .Y(n859) );
  NAND2X1 U1270 ( .A(\mem<18><1> ), .B(n25), .Y(n1532) );
  OAI21X1 U1271 ( .A(n145), .B(n1278), .C(n1532), .Y(n860) );
  NAND2X1 U1272 ( .A(\mem<18><2> ), .B(n25), .Y(n1533) );
  OAI21X1 U1273 ( .A(n145), .B(n1280), .C(n1533), .Y(n861) );
  NAND2X1 U1274 ( .A(\mem<18><3> ), .B(n25), .Y(n1534) );
  OAI21X1 U1275 ( .A(n145), .B(n1282), .C(n1534), .Y(n862) );
  NAND2X1 U1276 ( .A(\mem<18><4> ), .B(n25), .Y(n1535) );
  OAI21X1 U1277 ( .A(n145), .B(n1284), .C(n1535), .Y(n863) );
  NAND2X1 U1278 ( .A(\mem<18><5> ), .B(n25), .Y(n1536) );
  OAI21X1 U1279 ( .A(n145), .B(n1286), .C(n1536), .Y(n864) );
  NAND2X1 U1280 ( .A(\mem<18><6> ), .B(n25), .Y(n1537) );
  OAI21X1 U1281 ( .A(n145), .B(n1288), .C(n1537), .Y(n865) );
  NAND2X1 U1282 ( .A(\mem<18><7> ), .B(n25), .Y(n1538) );
  OAI21X1 U1283 ( .A(n145), .B(n1290), .C(n1538), .Y(n866) );
  NAND2X1 U1284 ( .A(\mem<18><8> ), .B(n25), .Y(n1539) );
  OAI21X1 U1285 ( .A(n145), .B(n1292), .C(n1539), .Y(n867) );
  NAND2X1 U1286 ( .A(\mem<18><9> ), .B(n25), .Y(n1540) );
  OAI21X1 U1287 ( .A(n145), .B(n1294), .C(n1540), .Y(n868) );
  NAND2X1 U1288 ( .A(\mem<18><10> ), .B(n25), .Y(n1541) );
  OAI21X1 U1289 ( .A(n145), .B(n1296), .C(n1541), .Y(n869) );
  NAND2X1 U1290 ( .A(\mem<18><11> ), .B(n25), .Y(n1542) );
  OAI21X1 U1291 ( .A(n145), .B(n1298), .C(n1542), .Y(n870) );
  NAND2X1 U1292 ( .A(\mem<18><12> ), .B(n25), .Y(n1543) );
  OAI21X1 U1293 ( .A(n145), .B(n1300), .C(n1543), .Y(n871) );
  NAND2X1 U1294 ( .A(\mem<18><13> ), .B(n25), .Y(n1544) );
  OAI21X1 U1295 ( .A(n145), .B(n1302), .C(n1544), .Y(n872) );
  NAND2X1 U1296 ( .A(\mem<18><14> ), .B(n25), .Y(n1545) );
  OAI21X1 U1297 ( .A(n145), .B(n1304), .C(n1545), .Y(n873) );
  NAND2X1 U1298 ( .A(\mem<18><15> ), .B(n25), .Y(n1546) );
  OAI21X1 U1299 ( .A(n145), .B(n1306), .C(n1546), .Y(n874) );
  NAND2X1 U1300 ( .A(\mem<17><0> ), .B(n27), .Y(n1547) );
  OAI21X1 U1301 ( .A(n147), .B(n1276), .C(n1547), .Y(n875) );
  NAND2X1 U1302 ( .A(\mem<17><1> ), .B(n27), .Y(n1548) );
  OAI21X1 U1303 ( .A(n147), .B(n1278), .C(n1548), .Y(n876) );
  NAND2X1 U1304 ( .A(\mem<17><2> ), .B(n27), .Y(n1549) );
  OAI21X1 U1305 ( .A(n147), .B(n1280), .C(n1549), .Y(n877) );
  NAND2X1 U1306 ( .A(\mem<17><3> ), .B(n27), .Y(n1550) );
  OAI21X1 U1307 ( .A(n147), .B(n1282), .C(n1550), .Y(n878) );
  NAND2X1 U1308 ( .A(\mem<17><4> ), .B(n27), .Y(n1551) );
  OAI21X1 U1309 ( .A(n147), .B(n1284), .C(n1551), .Y(n879) );
  NAND2X1 U1310 ( .A(\mem<17><5> ), .B(n27), .Y(n1552) );
  OAI21X1 U1311 ( .A(n147), .B(n1286), .C(n1552), .Y(n880) );
  NAND2X1 U1312 ( .A(\mem<17><6> ), .B(n27), .Y(n1553) );
  OAI21X1 U1313 ( .A(n147), .B(n1288), .C(n1553), .Y(n881) );
  NAND2X1 U1314 ( .A(\mem<17><7> ), .B(n27), .Y(n1554) );
  OAI21X1 U1315 ( .A(n147), .B(n1290), .C(n1554), .Y(n882) );
  NAND2X1 U1316 ( .A(\mem<17><8> ), .B(n27), .Y(n1555) );
  OAI21X1 U1317 ( .A(n147), .B(n1292), .C(n1555), .Y(n883) );
  NAND2X1 U1318 ( .A(\mem<17><9> ), .B(n27), .Y(n1556) );
  OAI21X1 U1319 ( .A(n147), .B(n1294), .C(n1556), .Y(n884) );
  NAND2X1 U1320 ( .A(\mem<17><10> ), .B(n27), .Y(n1557) );
  OAI21X1 U1321 ( .A(n147), .B(n1296), .C(n1557), .Y(n885) );
  NAND2X1 U1322 ( .A(\mem<17><11> ), .B(n27), .Y(n1558) );
  OAI21X1 U1323 ( .A(n147), .B(n1298), .C(n1558), .Y(n886) );
  NAND2X1 U1324 ( .A(\mem<17><12> ), .B(n27), .Y(n1559) );
  OAI21X1 U1325 ( .A(n147), .B(n1300), .C(n1559), .Y(n887) );
  NAND2X1 U1326 ( .A(\mem<17><13> ), .B(n27), .Y(n1560) );
  OAI21X1 U1327 ( .A(n147), .B(n1302), .C(n1560), .Y(n888) );
  NAND2X1 U1328 ( .A(\mem<17><14> ), .B(n27), .Y(n1561) );
  OAI21X1 U1329 ( .A(n147), .B(n1304), .C(n1561), .Y(n889) );
  NAND2X1 U1330 ( .A(\mem<17><15> ), .B(n27), .Y(n1562) );
  OAI21X1 U1331 ( .A(n147), .B(n1306), .C(n1562), .Y(n890) );
  NAND2X1 U1332 ( .A(\mem<16><0> ), .B(n29), .Y(n1563) );
  OAI21X1 U1333 ( .A(n1253), .B(n1276), .C(n1563), .Y(n891) );
  NAND2X1 U1334 ( .A(\mem<16><1> ), .B(n29), .Y(n1564) );
  OAI21X1 U1335 ( .A(n1253), .B(n1278), .C(n1564), .Y(n892) );
  NAND2X1 U1336 ( .A(\mem<16><2> ), .B(n29), .Y(n1565) );
  OAI21X1 U1337 ( .A(n1253), .B(n1280), .C(n1565), .Y(n893) );
  NAND2X1 U1338 ( .A(\mem<16><3> ), .B(n29), .Y(n1566) );
  OAI21X1 U1339 ( .A(n1253), .B(n1282), .C(n1566), .Y(n894) );
  NAND2X1 U1340 ( .A(\mem<16><4> ), .B(n29), .Y(n1567) );
  OAI21X1 U1341 ( .A(n1253), .B(n1284), .C(n1567), .Y(n895) );
  NAND2X1 U1342 ( .A(\mem<16><5> ), .B(n29), .Y(n1568) );
  OAI21X1 U1343 ( .A(n1253), .B(n1286), .C(n1568), .Y(n896) );
  NAND2X1 U1344 ( .A(\mem<16><6> ), .B(n29), .Y(n1569) );
  OAI21X1 U1345 ( .A(n1253), .B(n1288), .C(n1569), .Y(n897) );
  NAND2X1 U1346 ( .A(\mem<16><7> ), .B(n29), .Y(n1570) );
  OAI21X1 U1347 ( .A(n1253), .B(n1290), .C(n1570), .Y(n898) );
  NAND2X1 U1348 ( .A(\mem<16><8> ), .B(n29), .Y(n1571) );
  OAI21X1 U1349 ( .A(n1253), .B(n1292), .C(n1571), .Y(n899) );
  NAND2X1 U1350 ( .A(\mem<16><9> ), .B(n29), .Y(n1572) );
  OAI21X1 U1351 ( .A(n1253), .B(n1294), .C(n1572), .Y(n900) );
  NAND2X1 U1352 ( .A(\mem<16><10> ), .B(n29), .Y(n1573) );
  OAI21X1 U1353 ( .A(n1253), .B(n1296), .C(n1573), .Y(n901) );
  NAND2X1 U1354 ( .A(\mem<16><11> ), .B(n29), .Y(n1574) );
  OAI21X1 U1355 ( .A(n1253), .B(n1298), .C(n1574), .Y(n902) );
  NAND2X1 U1356 ( .A(\mem<16><12> ), .B(n29), .Y(n1575) );
  OAI21X1 U1357 ( .A(n1253), .B(n1300), .C(n1575), .Y(n903) );
  NAND2X1 U1358 ( .A(\mem<16><13> ), .B(n29), .Y(n1576) );
  OAI21X1 U1359 ( .A(n1253), .B(n1302), .C(n1576), .Y(n904) );
  NAND2X1 U1360 ( .A(\mem<16><14> ), .B(n29), .Y(n1577) );
  OAI21X1 U1361 ( .A(n1253), .B(n1304), .C(n1577), .Y(n905) );
  NAND2X1 U1362 ( .A(\mem<16><15> ), .B(n29), .Y(n1578) );
  OAI21X1 U1363 ( .A(n1253), .B(n1306), .C(n1578), .Y(n906) );
  NAND3X1 U1364 ( .A(n1187), .B(n214), .C(n1315), .Y(n1579) );
  NAND2X1 U1365 ( .A(\mem<15><0> ), .B(n31), .Y(n1580) );
  OAI21X1 U1366 ( .A(n149), .B(n1276), .C(n1580), .Y(n907) );
  NAND2X1 U1367 ( .A(\mem<15><1> ), .B(n31), .Y(n1581) );
  OAI21X1 U1368 ( .A(n149), .B(n1278), .C(n1581), .Y(n908) );
  NAND2X1 U1369 ( .A(\mem<15><2> ), .B(n31), .Y(n1582) );
  OAI21X1 U1370 ( .A(n149), .B(n1280), .C(n1582), .Y(n909) );
  NAND2X1 U1371 ( .A(\mem<15><3> ), .B(n31), .Y(n1583) );
  OAI21X1 U1372 ( .A(n149), .B(n1282), .C(n1583), .Y(n910) );
  NAND2X1 U1373 ( .A(\mem<15><4> ), .B(n31), .Y(n1584) );
  OAI21X1 U1374 ( .A(n149), .B(n1284), .C(n1584), .Y(n911) );
  NAND2X1 U1375 ( .A(\mem<15><5> ), .B(n31), .Y(n1585) );
  OAI21X1 U1376 ( .A(n149), .B(n1286), .C(n1585), .Y(n912) );
  NAND2X1 U1377 ( .A(\mem<15><6> ), .B(n31), .Y(n1586) );
  OAI21X1 U1378 ( .A(n149), .B(n1288), .C(n1586), .Y(n913) );
  NAND2X1 U1379 ( .A(\mem<15><7> ), .B(n31), .Y(n1587) );
  OAI21X1 U1380 ( .A(n149), .B(n1290), .C(n1587), .Y(n914) );
  NAND2X1 U1381 ( .A(\mem<15><8> ), .B(n31), .Y(n1588) );
  OAI21X1 U1382 ( .A(n149), .B(n1292), .C(n1588), .Y(n915) );
  NAND2X1 U1383 ( .A(\mem<15><9> ), .B(n31), .Y(n1589) );
  OAI21X1 U1384 ( .A(n149), .B(n1294), .C(n1589), .Y(n916) );
  NAND2X1 U1385 ( .A(\mem<15><10> ), .B(n31), .Y(n1590) );
  OAI21X1 U1386 ( .A(n149), .B(n1296), .C(n1590), .Y(n917) );
  NAND2X1 U1387 ( .A(\mem<15><11> ), .B(n31), .Y(n1591) );
  OAI21X1 U1388 ( .A(n149), .B(n1298), .C(n1591), .Y(n918) );
  NAND2X1 U1389 ( .A(\mem<15><12> ), .B(n31), .Y(n1592) );
  OAI21X1 U1390 ( .A(n149), .B(n1300), .C(n1592), .Y(n919) );
  NAND2X1 U1391 ( .A(\mem<15><13> ), .B(n31), .Y(n1593) );
  OAI21X1 U1392 ( .A(n149), .B(n1302), .C(n1593), .Y(n920) );
  NAND2X1 U1393 ( .A(\mem<15><14> ), .B(n31), .Y(n1594) );
  OAI21X1 U1394 ( .A(n149), .B(n1304), .C(n1594), .Y(n921) );
  NAND2X1 U1395 ( .A(\mem<15><15> ), .B(n31), .Y(n1595) );
  OAI21X1 U1396 ( .A(n149), .B(n1306), .C(n1595), .Y(n922) );
  NAND2X1 U1397 ( .A(\mem<14><0> ), .B(n33), .Y(n1596) );
  OAI21X1 U1398 ( .A(n151), .B(n1276), .C(n1596), .Y(n923) );
  NAND2X1 U1399 ( .A(\mem<14><1> ), .B(n33), .Y(n1597) );
  OAI21X1 U1400 ( .A(n151), .B(n1278), .C(n1597), .Y(n924) );
  NAND2X1 U1401 ( .A(\mem<14><2> ), .B(n33), .Y(n1598) );
  OAI21X1 U1402 ( .A(n151), .B(n1280), .C(n1598), .Y(n925) );
  NAND2X1 U1403 ( .A(\mem<14><3> ), .B(n33), .Y(n1599) );
  OAI21X1 U1404 ( .A(n151), .B(n1282), .C(n1599), .Y(n926) );
  NAND2X1 U1405 ( .A(\mem<14><4> ), .B(n33), .Y(n1600) );
  OAI21X1 U1406 ( .A(n151), .B(n1284), .C(n1600), .Y(n927) );
  NAND2X1 U1407 ( .A(\mem<14><5> ), .B(n33), .Y(n1601) );
  OAI21X1 U1408 ( .A(n151), .B(n1286), .C(n1601), .Y(n928) );
  NAND2X1 U1409 ( .A(\mem<14><6> ), .B(n33), .Y(n1602) );
  OAI21X1 U1410 ( .A(n151), .B(n1288), .C(n1602), .Y(n929) );
  NAND2X1 U1411 ( .A(\mem<14><7> ), .B(n33), .Y(n1603) );
  OAI21X1 U1412 ( .A(n151), .B(n1290), .C(n1603), .Y(n930) );
  NAND2X1 U1413 ( .A(\mem<14><8> ), .B(n33), .Y(n1604) );
  OAI21X1 U1414 ( .A(n151), .B(n1292), .C(n1604), .Y(n931) );
  NAND2X1 U1415 ( .A(\mem<14><9> ), .B(n33), .Y(n1605) );
  OAI21X1 U1416 ( .A(n151), .B(n1294), .C(n1605), .Y(n932) );
  NAND2X1 U1417 ( .A(\mem<14><10> ), .B(n33), .Y(n1606) );
  OAI21X1 U1418 ( .A(n151), .B(n1296), .C(n1606), .Y(n933) );
  NAND2X1 U1419 ( .A(\mem<14><11> ), .B(n33), .Y(n1607) );
  OAI21X1 U1420 ( .A(n151), .B(n1298), .C(n1607), .Y(n934) );
  NAND2X1 U1421 ( .A(\mem<14><12> ), .B(n33), .Y(n1608) );
  OAI21X1 U1422 ( .A(n151), .B(n1300), .C(n1608), .Y(n935) );
  NAND2X1 U1423 ( .A(\mem<14><13> ), .B(n33), .Y(n1609) );
  OAI21X1 U1424 ( .A(n151), .B(n1302), .C(n1609), .Y(n936) );
  NAND2X1 U1425 ( .A(\mem<14><14> ), .B(n33), .Y(n1610) );
  OAI21X1 U1426 ( .A(n151), .B(n1304), .C(n1610), .Y(n937) );
  NAND2X1 U1427 ( .A(\mem<14><15> ), .B(n33), .Y(n1611) );
  OAI21X1 U1428 ( .A(n151), .B(n1306), .C(n1611), .Y(n938) );
  NAND2X1 U1429 ( .A(\mem<13><0> ), .B(n35), .Y(n1612) );
  OAI21X1 U1430 ( .A(n153), .B(n1276), .C(n1612), .Y(n939) );
  NAND2X1 U1431 ( .A(\mem<13><1> ), .B(n35), .Y(n1613) );
  OAI21X1 U1432 ( .A(n153), .B(n1278), .C(n1613), .Y(n940) );
  NAND2X1 U1433 ( .A(\mem<13><2> ), .B(n35), .Y(n1614) );
  OAI21X1 U1434 ( .A(n153), .B(n1280), .C(n1614), .Y(n941) );
  NAND2X1 U1435 ( .A(\mem<13><3> ), .B(n35), .Y(n1615) );
  OAI21X1 U1436 ( .A(n153), .B(n1282), .C(n1615), .Y(n942) );
  NAND2X1 U1437 ( .A(\mem<13><4> ), .B(n35), .Y(n1616) );
  OAI21X1 U1438 ( .A(n153), .B(n1284), .C(n1616), .Y(n943) );
  NAND2X1 U1439 ( .A(\mem<13><5> ), .B(n35), .Y(n1617) );
  OAI21X1 U1440 ( .A(n153), .B(n1286), .C(n1617), .Y(n944) );
  NAND2X1 U1441 ( .A(\mem<13><6> ), .B(n35), .Y(n1618) );
  OAI21X1 U1442 ( .A(n153), .B(n1288), .C(n1618), .Y(n945) );
  NAND2X1 U1443 ( .A(\mem<13><7> ), .B(n35), .Y(n1619) );
  OAI21X1 U1444 ( .A(n153), .B(n1290), .C(n1619), .Y(n946) );
  NAND2X1 U1445 ( .A(\mem<13><8> ), .B(n35), .Y(n1620) );
  OAI21X1 U1446 ( .A(n153), .B(n1292), .C(n1620), .Y(n947) );
  NAND2X1 U1447 ( .A(\mem<13><9> ), .B(n35), .Y(n1621) );
  OAI21X1 U1448 ( .A(n153), .B(n1294), .C(n1621), .Y(n948) );
  NAND2X1 U1449 ( .A(\mem<13><10> ), .B(n35), .Y(n1622) );
  OAI21X1 U1450 ( .A(n153), .B(n1296), .C(n1622), .Y(n949) );
  NAND2X1 U1451 ( .A(\mem<13><11> ), .B(n35), .Y(n1623) );
  OAI21X1 U1452 ( .A(n153), .B(n1298), .C(n1623), .Y(n950) );
  NAND2X1 U1453 ( .A(\mem<13><12> ), .B(n35), .Y(n1624) );
  OAI21X1 U1454 ( .A(n153), .B(n1300), .C(n1624), .Y(n951) );
  NAND2X1 U1455 ( .A(\mem<13><13> ), .B(n35), .Y(n1625) );
  OAI21X1 U1456 ( .A(n153), .B(n1302), .C(n1625), .Y(n952) );
  NAND2X1 U1457 ( .A(\mem<13><14> ), .B(n35), .Y(n1626) );
  OAI21X1 U1458 ( .A(n153), .B(n1304), .C(n1626), .Y(n953) );
  NAND2X1 U1459 ( .A(\mem<13><15> ), .B(n35), .Y(n1627) );
  OAI21X1 U1460 ( .A(n153), .B(n1306), .C(n1627), .Y(n954) );
  NAND2X1 U1461 ( .A(\mem<12><0> ), .B(n37), .Y(n1628) );
  OAI21X1 U1462 ( .A(n155), .B(n1276), .C(n1628), .Y(n955) );
  NAND2X1 U1463 ( .A(\mem<12><1> ), .B(n37), .Y(n1629) );
  OAI21X1 U1464 ( .A(n155), .B(n1278), .C(n1629), .Y(n956) );
  NAND2X1 U1465 ( .A(\mem<12><2> ), .B(n37), .Y(n1630) );
  OAI21X1 U1466 ( .A(n155), .B(n1280), .C(n1630), .Y(n957) );
  NAND2X1 U1467 ( .A(\mem<12><3> ), .B(n37), .Y(n1631) );
  OAI21X1 U1468 ( .A(n155), .B(n1282), .C(n1631), .Y(n958) );
  NAND2X1 U1469 ( .A(\mem<12><4> ), .B(n37), .Y(n1632) );
  OAI21X1 U1470 ( .A(n155), .B(n1284), .C(n1632), .Y(n959) );
  NAND2X1 U1471 ( .A(\mem<12><5> ), .B(n37), .Y(n1633) );
  OAI21X1 U1472 ( .A(n155), .B(n1286), .C(n1633), .Y(n960) );
  NAND2X1 U1473 ( .A(\mem<12><6> ), .B(n37), .Y(n1634) );
  OAI21X1 U1474 ( .A(n155), .B(n1288), .C(n1634), .Y(n961) );
  NAND2X1 U1475 ( .A(\mem<12><7> ), .B(n37), .Y(n1635) );
  OAI21X1 U1476 ( .A(n155), .B(n1290), .C(n1635), .Y(n962) );
  NAND2X1 U1477 ( .A(\mem<12><8> ), .B(n37), .Y(n1636) );
  OAI21X1 U1478 ( .A(n155), .B(n1292), .C(n1636), .Y(n963) );
  NAND2X1 U1479 ( .A(\mem<12><9> ), .B(n37), .Y(n1637) );
  OAI21X1 U1480 ( .A(n155), .B(n1294), .C(n1637), .Y(n964) );
  NAND2X1 U1481 ( .A(\mem<12><10> ), .B(n37), .Y(n1638) );
  OAI21X1 U1482 ( .A(n155), .B(n1296), .C(n1638), .Y(n965) );
  NAND2X1 U1483 ( .A(\mem<12><11> ), .B(n37), .Y(n1639) );
  OAI21X1 U1484 ( .A(n155), .B(n1298), .C(n1639), .Y(n966) );
  NAND2X1 U1485 ( .A(\mem<12><12> ), .B(n37), .Y(n1640) );
  OAI21X1 U1486 ( .A(n155), .B(n1300), .C(n1640), .Y(n967) );
  NAND2X1 U1487 ( .A(\mem<12><13> ), .B(n37), .Y(n1641) );
  OAI21X1 U1488 ( .A(n155), .B(n1302), .C(n1641), .Y(n968) );
  NAND2X1 U1489 ( .A(\mem<12><14> ), .B(n37), .Y(n1642) );
  OAI21X1 U1490 ( .A(n155), .B(n1304), .C(n1642), .Y(n969) );
  NAND2X1 U1491 ( .A(\mem<12><15> ), .B(n37), .Y(n1643) );
  OAI21X1 U1492 ( .A(n155), .B(n1306), .C(n1643), .Y(n970) );
  NAND2X1 U1493 ( .A(\mem<11><0> ), .B(n39), .Y(n1644) );
  OAI21X1 U1494 ( .A(n157), .B(n1276), .C(n1644), .Y(n971) );
  NAND2X1 U1495 ( .A(\mem<11><1> ), .B(n39), .Y(n1645) );
  OAI21X1 U1496 ( .A(n157), .B(n1277), .C(n1645), .Y(n972) );
  NAND2X1 U1497 ( .A(\mem<11><2> ), .B(n39), .Y(n1646) );
  OAI21X1 U1498 ( .A(n157), .B(n1279), .C(n1646), .Y(n973) );
  NAND2X1 U1499 ( .A(\mem<11><3> ), .B(n39), .Y(n1647) );
  OAI21X1 U1500 ( .A(n157), .B(n1281), .C(n1647), .Y(n974) );
  NAND2X1 U1501 ( .A(\mem<11><4> ), .B(n39), .Y(n1648) );
  OAI21X1 U1502 ( .A(n157), .B(n1283), .C(n1648), .Y(n975) );
  NAND2X1 U1503 ( .A(\mem<11><5> ), .B(n39), .Y(n1649) );
  OAI21X1 U1504 ( .A(n157), .B(n1285), .C(n1649), .Y(n976) );
  NAND2X1 U1505 ( .A(\mem<11><6> ), .B(n39), .Y(n1650) );
  OAI21X1 U1506 ( .A(n157), .B(n1287), .C(n1650), .Y(n977) );
  NAND2X1 U1507 ( .A(\mem<11><7> ), .B(n39), .Y(n1651) );
  OAI21X1 U1508 ( .A(n157), .B(n1289), .C(n1651), .Y(n978) );
  NAND2X1 U1509 ( .A(\mem<11><8> ), .B(n39), .Y(n1652) );
  OAI21X1 U1510 ( .A(n157), .B(n1291), .C(n1652), .Y(n979) );
  NAND2X1 U1511 ( .A(\mem<11><9> ), .B(n39), .Y(n1653) );
  OAI21X1 U1512 ( .A(n157), .B(n1293), .C(n1653), .Y(n980) );
  NAND2X1 U1513 ( .A(\mem<11><10> ), .B(n39), .Y(n1654) );
  OAI21X1 U1514 ( .A(n157), .B(n1295), .C(n1654), .Y(n981) );
  NAND2X1 U1515 ( .A(\mem<11><11> ), .B(n39), .Y(n1655) );
  OAI21X1 U1516 ( .A(n157), .B(n1297), .C(n1655), .Y(n982) );
  NAND2X1 U1517 ( .A(\mem<11><12> ), .B(n39), .Y(n1656) );
  OAI21X1 U1518 ( .A(n157), .B(n1299), .C(n1656), .Y(n983) );
  NAND2X1 U1519 ( .A(\mem<11><13> ), .B(n39), .Y(n1657) );
  OAI21X1 U1520 ( .A(n157), .B(n1301), .C(n1657), .Y(n984) );
  NAND2X1 U1521 ( .A(\mem<11><14> ), .B(n39), .Y(n1658) );
  OAI21X1 U1522 ( .A(n157), .B(n1303), .C(n1658), .Y(n985) );
  NAND2X1 U1523 ( .A(\mem<11><15> ), .B(n39), .Y(n1659) );
  OAI21X1 U1524 ( .A(n157), .B(n1305), .C(n1659), .Y(n986) );
  NAND2X1 U1525 ( .A(\mem<10><0> ), .B(n41), .Y(n1660) );
  OAI21X1 U1526 ( .A(n159), .B(n1276), .C(n1660), .Y(n987) );
  NAND2X1 U1527 ( .A(\mem<10><1> ), .B(n41), .Y(n1661) );
  OAI21X1 U1528 ( .A(n159), .B(n1277), .C(n1661), .Y(n988) );
  NAND2X1 U1529 ( .A(\mem<10><2> ), .B(n41), .Y(n1662) );
  OAI21X1 U1530 ( .A(n159), .B(n1279), .C(n1662), .Y(n989) );
  NAND2X1 U1531 ( .A(\mem<10><3> ), .B(n41), .Y(n1663) );
  OAI21X1 U1532 ( .A(n159), .B(n1281), .C(n1663), .Y(n990) );
  NAND2X1 U1533 ( .A(\mem<10><4> ), .B(n41), .Y(n1664) );
  OAI21X1 U1534 ( .A(n159), .B(n1283), .C(n1664), .Y(n991) );
  NAND2X1 U1535 ( .A(\mem<10><5> ), .B(n41), .Y(n1665) );
  OAI21X1 U1536 ( .A(n159), .B(n1285), .C(n1665), .Y(n992) );
  NAND2X1 U1537 ( .A(\mem<10><6> ), .B(n41), .Y(n1666) );
  OAI21X1 U1538 ( .A(n159), .B(n1287), .C(n1666), .Y(n993) );
  NAND2X1 U1539 ( .A(\mem<10><7> ), .B(n41), .Y(n1667) );
  OAI21X1 U1540 ( .A(n159), .B(n1289), .C(n1667), .Y(n994) );
  NAND2X1 U1541 ( .A(\mem<10><8> ), .B(n41), .Y(n1668) );
  OAI21X1 U1542 ( .A(n159), .B(n1291), .C(n1668), .Y(n995) );
  NAND2X1 U1543 ( .A(\mem<10><9> ), .B(n41), .Y(n1669) );
  OAI21X1 U1544 ( .A(n159), .B(n1293), .C(n1669), .Y(n996) );
  NAND2X1 U1545 ( .A(\mem<10><10> ), .B(n41), .Y(n1670) );
  OAI21X1 U1546 ( .A(n159), .B(n1295), .C(n1670), .Y(n997) );
  NAND2X1 U1547 ( .A(\mem<10><11> ), .B(n41), .Y(n1671) );
  OAI21X1 U1548 ( .A(n159), .B(n1297), .C(n1671), .Y(n998) );
  NAND2X1 U1549 ( .A(\mem<10><12> ), .B(n41), .Y(n1672) );
  OAI21X1 U1550 ( .A(n159), .B(n1299), .C(n1672), .Y(n999) );
  NAND2X1 U1551 ( .A(\mem<10><13> ), .B(n41), .Y(n1673) );
  OAI21X1 U1552 ( .A(n159), .B(n1301), .C(n1673), .Y(n1000) );
  NAND2X1 U1553 ( .A(\mem<10><14> ), .B(n41), .Y(n1674) );
  OAI21X1 U1554 ( .A(n159), .B(n1303), .C(n1674), .Y(n1001) );
  NAND2X1 U1555 ( .A(\mem<10><15> ), .B(n41), .Y(n1675) );
  OAI21X1 U1556 ( .A(n159), .B(n1305), .C(n1675), .Y(n1002) );
  NAND2X1 U1557 ( .A(\mem<9><0> ), .B(n43), .Y(n1676) );
  OAI21X1 U1558 ( .A(n161), .B(n1276), .C(n1676), .Y(n1003) );
  NAND2X1 U1559 ( .A(\mem<9><1> ), .B(n43), .Y(n1677) );
  OAI21X1 U1560 ( .A(n161), .B(n1277), .C(n1677), .Y(n1004) );
  NAND2X1 U1561 ( .A(\mem<9><2> ), .B(n43), .Y(n1678) );
  OAI21X1 U1562 ( .A(n161), .B(n1279), .C(n1678), .Y(n1005) );
  NAND2X1 U1563 ( .A(\mem<9><3> ), .B(n43), .Y(n1679) );
  OAI21X1 U1564 ( .A(n161), .B(n1281), .C(n1679), .Y(n1006) );
  NAND2X1 U1565 ( .A(\mem<9><4> ), .B(n43), .Y(n1680) );
  OAI21X1 U1566 ( .A(n161), .B(n1283), .C(n1680), .Y(n1007) );
  NAND2X1 U1567 ( .A(\mem<9><5> ), .B(n43), .Y(n1681) );
  OAI21X1 U1568 ( .A(n161), .B(n1285), .C(n1681), .Y(n1008) );
  NAND2X1 U1569 ( .A(\mem<9><6> ), .B(n43), .Y(n1682) );
  OAI21X1 U1570 ( .A(n161), .B(n1287), .C(n1682), .Y(n1009) );
  NAND2X1 U1571 ( .A(\mem<9><7> ), .B(n43), .Y(n1683) );
  OAI21X1 U1572 ( .A(n161), .B(n1289), .C(n1683), .Y(n1010) );
  NAND2X1 U1573 ( .A(\mem<9><8> ), .B(n43), .Y(n1684) );
  OAI21X1 U1574 ( .A(n161), .B(n1291), .C(n1684), .Y(n1011) );
  NAND2X1 U1575 ( .A(\mem<9><9> ), .B(n43), .Y(n1685) );
  OAI21X1 U1576 ( .A(n161), .B(n1293), .C(n1685), .Y(n1012) );
  NAND2X1 U1577 ( .A(\mem<9><10> ), .B(n43), .Y(n1686) );
  OAI21X1 U1578 ( .A(n161), .B(n1295), .C(n1686), .Y(n1013) );
  NAND2X1 U1579 ( .A(\mem<9><11> ), .B(n43), .Y(n1687) );
  OAI21X1 U1580 ( .A(n161), .B(n1297), .C(n1687), .Y(n1014) );
  NAND2X1 U1581 ( .A(\mem<9><12> ), .B(n43), .Y(n1688) );
  OAI21X1 U1582 ( .A(n161), .B(n1299), .C(n1688), .Y(n1015) );
  NAND2X1 U1583 ( .A(\mem<9><13> ), .B(n43), .Y(n1689) );
  OAI21X1 U1584 ( .A(n161), .B(n1301), .C(n1689), .Y(n1016) );
  NAND2X1 U1585 ( .A(\mem<9><14> ), .B(n43), .Y(n1690) );
  OAI21X1 U1586 ( .A(n161), .B(n1303), .C(n1690), .Y(n1017) );
  NAND2X1 U1587 ( .A(\mem<9><15> ), .B(n43), .Y(n1691) );
  OAI21X1 U1588 ( .A(n161), .B(n1305), .C(n1691), .Y(n1018) );
  NAND2X1 U1589 ( .A(\mem<8><0> ), .B(n102), .Y(n1693) );
  OAI21X1 U1590 ( .A(n1254), .B(n1276), .C(n1693), .Y(n1019) );
  NAND2X1 U1591 ( .A(\mem<8><1> ), .B(n102), .Y(n1694) );
  OAI21X1 U1592 ( .A(n1254), .B(n1277), .C(n1694), .Y(n1020) );
  NAND2X1 U1593 ( .A(\mem<8><2> ), .B(n102), .Y(n1695) );
  OAI21X1 U1594 ( .A(n1254), .B(n1279), .C(n1695), .Y(n1021) );
  NAND2X1 U1595 ( .A(\mem<8><3> ), .B(n102), .Y(n1696) );
  OAI21X1 U1596 ( .A(n1254), .B(n1281), .C(n1696), .Y(n1022) );
  NAND2X1 U1597 ( .A(\mem<8><4> ), .B(n102), .Y(n1697) );
  OAI21X1 U1598 ( .A(n1254), .B(n1283), .C(n1697), .Y(n1023) );
  NAND2X1 U1599 ( .A(\mem<8><5> ), .B(n102), .Y(n1698) );
  OAI21X1 U1600 ( .A(n1254), .B(n1285), .C(n1698), .Y(n1024) );
  NAND2X1 U1601 ( .A(\mem<8><6> ), .B(n102), .Y(n1699) );
  OAI21X1 U1602 ( .A(n1254), .B(n1287), .C(n1699), .Y(n1025) );
  NAND2X1 U1603 ( .A(\mem<8><7> ), .B(n102), .Y(n1700) );
  OAI21X1 U1604 ( .A(n1254), .B(n1289), .C(n1700), .Y(n1026) );
  NAND2X1 U1605 ( .A(\mem<8><8> ), .B(n102), .Y(n1701) );
  OAI21X1 U1606 ( .A(n1254), .B(n1291), .C(n1701), .Y(n1027) );
  NAND2X1 U1607 ( .A(\mem<8><9> ), .B(n102), .Y(n1702) );
  OAI21X1 U1608 ( .A(n1254), .B(n1293), .C(n1702), .Y(n1028) );
  NAND2X1 U1609 ( .A(\mem<8><10> ), .B(n102), .Y(n1703) );
  OAI21X1 U1610 ( .A(n1254), .B(n1295), .C(n1703), .Y(n1029) );
  NAND2X1 U1611 ( .A(\mem<8><11> ), .B(n102), .Y(n1704) );
  OAI21X1 U1612 ( .A(n1254), .B(n1297), .C(n1704), .Y(n1030) );
  NAND2X1 U1613 ( .A(\mem<8><12> ), .B(n102), .Y(n1705) );
  OAI21X1 U1614 ( .A(n1254), .B(n1299), .C(n1705), .Y(n1031) );
  NAND2X1 U1615 ( .A(\mem<8><13> ), .B(n102), .Y(n1706) );
  OAI21X1 U1616 ( .A(n1254), .B(n1301), .C(n1706), .Y(n1032) );
  NAND2X1 U1617 ( .A(\mem<8><14> ), .B(n102), .Y(n1707) );
  OAI21X1 U1618 ( .A(n1254), .B(n1303), .C(n1707), .Y(n1033) );
  NAND2X1 U1619 ( .A(\mem<8><15> ), .B(n102), .Y(n1708) );
  OAI21X1 U1620 ( .A(n1254), .B(n1305), .C(n1708), .Y(n1034) );
  NAND3X1 U1621 ( .A(n1313), .B(n214), .C(n1315), .Y(n1709) );
  NAND2X1 U1622 ( .A(\mem<7><0> ), .B(n1255), .Y(n1710) );
  OAI21X1 U1623 ( .A(n163), .B(n1275), .C(n1710), .Y(n1035) );
  NAND2X1 U1624 ( .A(\mem<7><1> ), .B(n19), .Y(n1711) );
  OAI21X1 U1625 ( .A(n163), .B(n1277), .C(n1711), .Y(n1036) );
  NAND2X1 U1626 ( .A(\mem<7><2> ), .B(n1256), .Y(n1712) );
  OAI21X1 U1627 ( .A(n163), .B(n1279), .C(n1712), .Y(n1037) );
  NAND2X1 U1628 ( .A(\mem<7><3> ), .B(n1255), .Y(n1713) );
  OAI21X1 U1629 ( .A(n163), .B(n1281), .C(n1713), .Y(n1038) );
  NAND2X1 U1630 ( .A(\mem<7><4> ), .B(n19), .Y(n1714) );
  OAI21X1 U1631 ( .A(n163), .B(n1283), .C(n1714), .Y(n1039) );
  NAND2X1 U1632 ( .A(\mem<7><5> ), .B(n1256), .Y(n1715) );
  OAI21X1 U1633 ( .A(n163), .B(n1285), .C(n1715), .Y(n1040) );
  NAND2X1 U1634 ( .A(\mem<7><6> ), .B(n1255), .Y(n1716) );
  OAI21X1 U1635 ( .A(n163), .B(n1287), .C(n1716), .Y(n1041) );
  NAND2X1 U1636 ( .A(\mem<7><7> ), .B(n19), .Y(n1717) );
  OAI21X1 U1637 ( .A(n163), .B(n1289), .C(n1717), .Y(n1042) );
  NAND2X1 U1638 ( .A(\mem<7><8> ), .B(n1256), .Y(n1718) );
  OAI21X1 U1639 ( .A(n163), .B(n1291), .C(n1718), .Y(n1043) );
  NAND2X1 U1640 ( .A(\mem<7><9> ), .B(n1255), .Y(n1719) );
  OAI21X1 U1641 ( .A(n163), .B(n1293), .C(n1719), .Y(n1044) );
  NAND2X1 U1642 ( .A(\mem<7><10> ), .B(n19), .Y(n1720) );
  OAI21X1 U1643 ( .A(n163), .B(n1295), .C(n1720), .Y(n1045) );
  NAND2X1 U1644 ( .A(\mem<7><11> ), .B(n1256), .Y(n1721) );
  OAI21X1 U1645 ( .A(n163), .B(n1297), .C(n1721), .Y(n1046) );
  NAND2X1 U1646 ( .A(\mem<7><12> ), .B(n1255), .Y(n1722) );
  OAI21X1 U1647 ( .A(n163), .B(n1299), .C(n1722), .Y(n1047) );
  NAND2X1 U1648 ( .A(\mem<7><13> ), .B(n19), .Y(n1723) );
  OAI21X1 U1649 ( .A(n163), .B(n1301), .C(n1723), .Y(n1048) );
  NAND2X1 U1650 ( .A(\mem<7><14> ), .B(n1256), .Y(n1724) );
  OAI21X1 U1651 ( .A(n163), .B(n1303), .C(n1724), .Y(n1049) );
  NAND2X1 U1652 ( .A(\mem<7><15> ), .B(n1255), .Y(n1725) );
  OAI21X1 U1653 ( .A(n163), .B(n1305), .C(n1725), .Y(n1050) );
  NAND2X1 U1654 ( .A(\mem<6><0> ), .B(n1257), .Y(n1726) );
  OAI21X1 U1655 ( .A(n165), .B(n1276), .C(n1726), .Y(n1051) );
  NAND2X1 U1656 ( .A(\mem<6><1> ), .B(n18), .Y(n1727) );
  OAI21X1 U1657 ( .A(n165), .B(n1277), .C(n1727), .Y(n1052) );
  NAND2X1 U1658 ( .A(\mem<6><2> ), .B(n1258), .Y(n1728) );
  OAI21X1 U1659 ( .A(n165), .B(n1279), .C(n1728), .Y(n1053) );
  NAND2X1 U1660 ( .A(\mem<6><3> ), .B(n1257), .Y(n1729) );
  OAI21X1 U1661 ( .A(n165), .B(n1281), .C(n1729), .Y(n1054) );
  NAND2X1 U1662 ( .A(\mem<6><4> ), .B(n18), .Y(n1730) );
  OAI21X1 U1663 ( .A(n165), .B(n1283), .C(n1730), .Y(n1055) );
  NAND2X1 U1664 ( .A(\mem<6><5> ), .B(n1258), .Y(n1731) );
  OAI21X1 U1665 ( .A(n165), .B(n1285), .C(n1731), .Y(n1056) );
  NAND2X1 U1666 ( .A(\mem<6><6> ), .B(n1257), .Y(n1732) );
  OAI21X1 U1667 ( .A(n165), .B(n1287), .C(n1732), .Y(n1057) );
  NAND2X1 U1668 ( .A(\mem<6><7> ), .B(n18), .Y(n1733) );
  OAI21X1 U1669 ( .A(n165), .B(n1289), .C(n1733), .Y(n1058) );
  NAND2X1 U1670 ( .A(\mem<6><8> ), .B(n1258), .Y(n1734) );
  OAI21X1 U1671 ( .A(n165), .B(n1291), .C(n1734), .Y(n1059) );
  NAND2X1 U1672 ( .A(\mem<6><9> ), .B(n1257), .Y(n1735) );
  OAI21X1 U1673 ( .A(n165), .B(n1293), .C(n1735), .Y(n1060) );
  NAND2X1 U1674 ( .A(\mem<6><10> ), .B(n18), .Y(n1736) );
  OAI21X1 U1675 ( .A(n165), .B(n1295), .C(n1736), .Y(n1061) );
  NAND2X1 U1676 ( .A(\mem<6><11> ), .B(n1258), .Y(n1737) );
  OAI21X1 U1677 ( .A(n165), .B(n1297), .C(n1737), .Y(n1062) );
  NAND2X1 U1678 ( .A(\mem<6><12> ), .B(n1257), .Y(n1738) );
  OAI21X1 U1679 ( .A(n165), .B(n1299), .C(n1738), .Y(n1063) );
  NAND2X1 U1680 ( .A(\mem<6><13> ), .B(n18), .Y(n1739) );
  OAI21X1 U1681 ( .A(n165), .B(n1301), .C(n1739), .Y(n1064) );
  NAND2X1 U1682 ( .A(\mem<6><14> ), .B(n1258), .Y(n1740) );
  OAI21X1 U1683 ( .A(n165), .B(n1303), .C(n1740), .Y(n1065) );
  NAND2X1 U1684 ( .A(\mem<6><15> ), .B(n1257), .Y(n1741) );
  OAI21X1 U1685 ( .A(n165), .B(n1305), .C(n1741), .Y(n1066) );
  NAND2X1 U1686 ( .A(\mem<5><0> ), .B(n1259), .Y(n1743) );
  OAI21X1 U1687 ( .A(n167), .B(n1275), .C(n1743), .Y(n1067) );
  NAND2X1 U1688 ( .A(\mem<5><1> ), .B(n17), .Y(n1744) );
  OAI21X1 U1689 ( .A(n167), .B(n1277), .C(n1744), .Y(n1068) );
  NAND2X1 U1690 ( .A(\mem<5><2> ), .B(n1260), .Y(n1745) );
  OAI21X1 U1691 ( .A(n167), .B(n1279), .C(n1745), .Y(n1069) );
  NAND2X1 U1692 ( .A(\mem<5><3> ), .B(n1259), .Y(n1746) );
  OAI21X1 U1693 ( .A(n167), .B(n1281), .C(n1746), .Y(n1070) );
  NAND2X1 U1694 ( .A(\mem<5><4> ), .B(n17), .Y(n1747) );
  OAI21X1 U1695 ( .A(n167), .B(n1283), .C(n1747), .Y(n1071) );
  NAND2X1 U1696 ( .A(\mem<5><5> ), .B(n1260), .Y(n1748) );
  OAI21X1 U1697 ( .A(n167), .B(n1285), .C(n1748), .Y(n1072) );
  NAND2X1 U1698 ( .A(\mem<5><6> ), .B(n1259), .Y(n1749) );
  OAI21X1 U1699 ( .A(n167), .B(n1287), .C(n1749), .Y(n1073) );
  NAND2X1 U1700 ( .A(\mem<5><7> ), .B(n17), .Y(n1750) );
  OAI21X1 U1701 ( .A(n167), .B(n1289), .C(n1750), .Y(n1074) );
  NAND2X1 U1702 ( .A(\mem<5><8> ), .B(n1260), .Y(n1751) );
  OAI21X1 U1703 ( .A(n167), .B(n1291), .C(n1751), .Y(n1075) );
  NAND2X1 U1704 ( .A(\mem<5><9> ), .B(n1259), .Y(n1752) );
  OAI21X1 U1705 ( .A(n167), .B(n1293), .C(n1752), .Y(n1076) );
  NAND2X1 U1706 ( .A(\mem<5><10> ), .B(n17), .Y(n1753) );
  OAI21X1 U1707 ( .A(n167), .B(n1295), .C(n1753), .Y(n1077) );
  NAND2X1 U1708 ( .A(\mem<5><11> ), .B(n1260), .Y(n1754) );
  OAI21X1 U1709 ( .A(n167), .B(n1297), .C(n1754), .Y(n1078) );
  NAND2X1 U1710 ( .A(\mem<5><12> ), .B(n1259), .Y(n1755) );
  OAI21X1 U1711 ( .A(n167), .B(n1299), .C(n1755), .Y(n1079) );
  NAND2X1 U1712 ( .A(\mem<5><13> ), .B(n17), .Y(n1756) );
  OAI21X1 U1713 ( .A(n167), .B(n1301), .C(n1756), .Y(n1080) );
  NAND2X1 U1714 ( .A(\mem<5><14> ), .B(n1260), .Y(n1757) );
  OAI21X1 U1715 ( .A(n167), .B(n1303), .C(n1757), .Y(n1081) );
  NAND2X1 U1716 ( .A(\mem<5><15> ), .B(n1259), .Y(n1758) );
  OAI21X1 U1717 ( .A(n167), .B(n1305), .C(n1758), .Y(n1082) );
  NAND2X1 U1718 ( .A(\mem<4><0> ), .B(n1261), .Y(n1760) );
  OAI21X1 U1719 ( .A(n169), .B(n1276), .C(n1760), .Y(n1083) );
  NAND2X1 U1720 ( .A(\mem<4><1> ), .B(n16), .Y(n1761) );
  OAI21X1 U1721 ( .A(n169), .B(n1277), .C(n1761), .Y(n1084) );
  NAND2X1 U1722 ( .A(\mem<4><2> ), .B(n1262), .Y(n1762) );
  OAI21X1 U1723 ( .A(n169), .B(n1279), .C(n1762), .Y(n1085) );
  NAND2X1 U1724 ( .A(\mem<4><3> ), .B(n1261), .Y(n1763) );
  OAI21X1 U1725 ( .A(n169), .B(n1281), .C(n1763), .Y(n1086) );
  NAND2X1 U1726 ( .A(\mem<4><4> ), .B(n16), .Y(n1764) );
  OAI21X1 U1727 ( .A(n169), .B(n1283), .C(n1764), .Y(n1087) );
  NAND2X1 U1728 ( .A(\mem<4><5> ), .B(n1262), .Y(n1765) );
  OAI21X1 U1729 ( .A(n169), .B(n1285), .C(n1765), .Y(n1088) );
  NAND2X1 U1730 ( .A(\mem<4><6> ), .B(n1261), .Y(n1766) );
  OAI21X1 U1731 ( .A(n169), .B(n1287), .C(n1766), .Y(n1089) );
  NAND2X1 U1732 ( .A(\mem<4><7> ), .B(n16), .Y(n1767) );
  OAI21X1 U1733 ( .A(n169), .B(n1289), .C(n1767), .Y(n1090) );
  NAND2X1 U1734 ( .A(\mem<4><8> ), .B(n1262), .Y(n1768) );
  OAI21X1 U1735 ( .A(n169), .B(n1291), .C(n1768), .Y(n1091) );
  NAND2X1 U1736 ( .A(\mem<4><9> ), .B(n1261), .Y(n1769) );
  OAI21X1 U1737 ( .A(n169), .B(n1293), .C(n1769), .Y(n1092) );
  NAND2X1 U1738 ( .A(\mem<4><10> ), .B(n16), .Y(n1770) );
  OAI21X1 U1739 ( .A(n169), .B(n1295), .C(n1770), .Y(n1093) );
  NAND2X1 U1740 ( .A(\mem<4><11> ), .B(n1262), .Y(n1771) );
  OAI21X1 U1741 ( .A(n169), .B(n1297), .C(n1771), .Y(n1094) );
  NAND2X1 U1742 ( .A(\mem<4><12> ), .B(n1261), .Y(n1772) );
  OAI21X1 U1743 ( .A(n169), .B(n1299), .C(n1772), .Y(n1095) );
  NAND2X1 U1744 ( .A(\mem<4><13> ), .B(n16), .Y(n1773) );
  OAI21X1 U1745 ( .A(n169), .B(n1301), .C(n1773), .Y(n1096) );
  NAND2X1 U1746 ( .A(\mem<4><14> ), .B(n1262), .Y(n1774) );
  OAI21X1 U1747 ( .A(n169), .B(n1303), .C(n1774), .Y(n1097) );
  NAND2X1 U1748 ( .A(\mem<4><15> ), .B(n1261), .Y(n1775) );
  OAI21X1 U1749 ( .A(n169), .B(n1305), .C(n1775), .Y(n1098) );
  NAND2X1 U1750 ( .A(\mem<3><0> ), .B(n1263), .Y(n1777) );
  OAI21X1 U1751 ( .A(n171), .B(n1275), .C(n1777), .Y(n1099) );
  NAND2X1 U1752 ( .A(\mem<3><1> ), .B(n15), .Y(n1778) );
  OAI21X1 U1753 ( .A(n171), .B(n1277), .C(n1778), .Y(n1100) );
  NAND2X1 U1754 ( .A(\mem<3><2> ), .B(n1264), .Y(n1779) );
  OAI21X1 U1755 ( .A(n171), .B(n1279), .C(n1779), .Y(n1101) );
  NAND2X1 U1756 ( .A(\mem<3><3> ), .B(n1263), .Y(n1780) );
  OAI21X1 U1757 ( .A(n171), .B(n1281), .C(n1780), .Y(n1102) );
  NAND2X1 U1758 ( .A(\mem<3><4> ), .B(n15), .Y(n1781) );
  OAI21X1 U1759 ( .A(n171), .B(n1283), .C(n1781), .Y(n1103) );
  NAND2X1 U1760 ( .A(\mem<3><5> ), .B(n1264), .Y(n1782) );
  OAI21X1 U1761 ( .A(n171), .B(n1285), .C(n1782), .Y(n1104) );
  NAND2X1 U1762 ( .A(\mem<3><6> ), .B(n1263), .Y(n1783) );
  OAI21X1 U1763 ( .A(n171), .B(n1287), .C(n1783), .Y(n1105) );
  NAND2X1 U1764 ( .A(\mem<3><7> ), .B(n15), .Y(n1784) );
  OAI21X1 U1765 ( .A(n171), .B(n1289), .C(n1784), .Y(n1106) );
  NAND2X1 U1766 ( .A(\mem<3><8> ), .B(n1264), .Y(n1785) );
  OAI21X1 U1767 ( .A(n171), .B(n1291), .C(n1785), .Y(n1107) );
  NAND2X1 U1768 ( .A(\mem<3><9> ), .B(n1263), .Y(n1786) );
  OAI21X1 U1769 ( .A(n171), .B(n1293), .C(n1786), .Y(n1108) );
  NAND2X1 U1770 ( .A(\mem<3><10> ), .B(n15), .Y(n1787) );
  OAI21X1 U1771 ( .A(n171), .B(n1295), .C(n1787), .Y(n1109) );
  NAND2X1 U1772 ( .A(\mem<3><11> ), .B(n1264), .Y(n1788) );
  OAI21X1 U1773 ( .A(n171), .B(n1297), .C(n1788), .Y(n1110) );
  NAND2X1 U1774 ( .A(\mem<3><12> ), .B(n1263), .Y(n1789) );
  OAI21X1 U1775 ( .A(n171), .B(n1299), .C(n1789), .Y(n1111) );
  NAND2X1 U1776 ( .A(\mem<3><13> ), .B(n15), .Y(n1790) );
  OAI21X1 U1777 ( .A(n171), .B(n1301), .C(n1790), .Y(n1112) );
  NAND2X1 U1778 ( .A(\mem<3><14> ), .B(n1264), .Y(n1791) );
  OAI21X1 U1779 ( .A(n171), .B(n1303), .C(n1791), .Y(n1113) );
  NAND2X1 U1780 ( .A(\mem<3><15> ), .B(n1263), .Y(n1792) );
  OAI21X1 U1781 ( .A(n171), .B(n1305), .C(n1792), .Y(n1114) );
  NAND2X1 U1782 ( .A(\mem<2><0> ), .B(n1265), .Y(n1794) );
  OAI21X1 U1783 ( .A(n173), .B(n1276), .C(n1794), .Y(n1115) );
  NAND2X1 U1784 ( .A(\mem<2><1> ), .B(n14), .Y(n1795) );
  OAI21X1 U1785 ( .A(n173), .B(n1277), .C(n1795), .Y(n1116) );
  NAND2X1 U1786 ( .A(\mem<2><2> ), .B(n1266), .Y(n1796) );
  OAI21X1 U1787 ( .A(n173), .B(n1279), .C(n1796), .Y(n1117) );
  NAND2X1 U1788 ( .A(\mem<2><3> ), .B(n1265), .Y(n1797) );
  OAI21X1 U1789 ( .A(n173), .B(n1281), .C(n1797), .Y(n1118) );
  NAND2X1 U1790 ( .A(\mem<2><4> ), .B(n14), .Y(n1798) );
  OAI21X1 U1791 ( .A(n173), .B(n1283), .C(n1798), .Y(n1119) );
  NAND2X1 U1792 ( .A(\mem<2><5> ), .B(n1266), .Y(n1799) );
  OAI21X1 U1793 ( .A(n173), .B(n1285), .C(n1799), .Y(n1120) );
  NAND2X1 U1794 ( .A(\mem<2><6> ), .B(n1265), .Y(n1800) );
  OAI21X1 U1795 ( .A(n173), .B(n1287), .C(n1800), .Y(n1121) );
  NAND2X1 U1796 ( .A(\mem<2><7> ), .B(n14), .Y(n1801) );
  OAI21X1 U1797 ( .A(n173), .B(n1289), .C(n1801), .Y(n1122) );
  NAND2X1 U1798 ( .A(\mem<2><8> ), .B(n1266), .Y(n1802) );
  OAI21X1 U1799 ( .A(n173), .B(n1291), .C(n1802), .Y(n1123) );
  NAND2X1 U1800 ( .A(\mem<2><9> ), .B(n1265), .Y(n1803) );
  OAI21X1 U1801 ( .A(n173), .B(n1293), .C(n1803), .Y(n1124) );
  NAND2X1 U1802 ( .A(\mem<2><10> ), .B(n14), .Y(n1804) );
  OAI21X1 U1803 ( .A(n173), .B(n1295), .C(n1804), .Y(n1125) );
  NAND2X1 U1804 ( .A(\mem<2><11> ), .B(n1266), .Y(n1805) );
  OAI21X1 U1805 ( .A(n173), .B(n1297), .C(n1805), .Y(n1126) );
  NAND2X1 U1806 ( .A(\mem<2><12> ), .B(n1265), .Y(n1806) );
  OAI21X1 U1807 ( .A(n173), .B(n1299), .C(n1806), .Y(n1127) );
  NAND2X1 U1808 ( .A(\mem<2><13> ), .B(n14), .Y(n1807) );
  OAI21X1 U1809 ( .A(n173), .B(n1301), .C(n1807), .Y(n1128) );
  NAND2X1 U1810 ( .A(\mem<2><14> ), .B(n1266), .Y(n1808) );
  OAI21X1 U1811 ( .A(n173), .B(n1303), .C(n1808), .Y(n1129) );
  NAND2X1 U1812 ( .A(\mem<2><15> ), .B(n1265), .Y(n1809) );
  OAI21X1 U1813 ( .A(n173), .B(n1305), .C(n1809), .Y(n1130) );
  NAND2X1 U1814 ( .A(\mem<1><0> ), .B(n1268), .Y(n1811) );
  OAI21X1 U1815 ( .A(n175), .B(n1275), .C(n1811), .Y(n1131) );
  NAND2X1 U1816 ( .A(\mem<1><1> ), .B(n13), .Y(n1812) );
  OAI21X1 U1817 ( .A(n175), .B(n1277), .C(n1812), .Y(n1132) );
  NAND2X1 U1818 ( .A(\mem<1><2> ), .B(n1268), .Y(n1813) );
  OAI21X1 U1819 ( .A(n175), .B(n1279), .C(n1813), .Y(n1133) );
  NAND2X1 U1820 ( .A(\mem<1><3> ), .B(n13), .Y(n1814) );
  OAI21X1 U1821 ( .A(n175), .B(n1281), .C(n1814), .Y(n1134) );
  NAND2X1 U1822 ( .A(\mem<1><4> ), .B(n1268), .Y(n1815) );
  OAI21X1 U1823 ( .A(n175), .B(n1283), .C(n1815), .Y(n1135) );
  NAND2X1 U1824 ( .A(\mem<1><5> ), .B(n13), .Y(n1816) );
  OAI21X1 U1825 ( .A(n175), .B(n1285), .C(n1816), .Y(n1136) );
  NAND2X1 U1826 ( .A(\mem<1><6> ), .B(n1268), .Y(n1817) );
  OAI21X1 U1827 ( .A(n175), .B(n1287), .C(n1817), .Y(n1137) );
  NAND2X1 U1828 ( .A(\mem<1><7> ), .B(n13), .Y(n1818) );
  OAI21X1 U1829 ( .A(n175), .B(n1289), .C(n1818), .Y(n1138) );
  NAND2X1 U1830 ( .A(\mem<1><8> ), .B(n1268), .Y(n1819) );
  OAI21X1 U1831 ( .A(n175), .B(n1291), .C(n1819), .Y(n1139) );
  NAND2X1 U1832 ( .A(\mem<1><9> ), .B(n13), .Y(n1820) );
  OAI21X1 U1833 ( .A(n175), .B(n1293), .C(n1820), .Y(n1140) );
  NAND2X1 U1834 ( .A(\mem<1><10> ), .B(n1267), .Y(n1821) );
  OAI21X1 U1835 ( .A(n175), .B(n1295), .C(n1821), .Y(n1141) );
  NAND2X1 U1836 ( .A(\mem<1><11> ), .B(n1267), .Y(n1822) );
  OAI21X1 U1837 ( .A(n175), .B(n1297), .C(n1822), .Y(n1142) );
  NAND2X1 U1838 ( .A(\mem<1><12> ), .B(n1267), .Y(n1823) );
  OAI21X1 U1839 ( .A(n175), .B(n1299), .C(n1823), .Y(n1143) );
  NAND2X1 U1840 ( .A(\mem<1><13> ), .B(n1267), .Y(n1824) );
  OAI21X1 U1841 ( .A(n175), .B(n1301), .C(n1824), .Y(n1144) );
  NAND2X1 U1842 ( .A(\mem<1><14> ), .B(n1267), .Y(n1825) );
  OAI21X1 U1843 ( .A(n175), .B(n1303), .C(n1825), .Y(n1145) );
  NAND2X1 U1844 ( .A(\mem<1><15> ), .B(n1267), .Y(n1826) );
  OAI21X1 U1845 ( .A(n175), .B(n1305), .C(n1826), .Y(n1146) );
  NAND2X1 U1846 ( .A(\mem<0><0> ), .B(n45), .Y(n1829) );
  OAI21X1 U1847 ( .A(n1269), .B(n1276), .C(n1829), .Y(n1147) );
  NAND2X1 U1848 ( .A(\mem<0><1> ), .B(n45), .Y(n1830) );
  OAI21X1 U1849 ( .A(n1269), .B(n1277), .C(n1830), .Y(n1148) );
  NAND2X1 U1850 ( .A(\mem<0><2> ), .B(n45), .Y(n1831) );
  OAI21X1 U1851 ( .A(n1269), .B(n1279), .C(n1831), .Y(n1149) );
  NAND2X1 U1852 ( .A(\mem<0><3> ), .B(n45), .Y(n1832) );
  OAI21X1 U1853 ( .A(n1269), .B(n1281), .C(n1832), .Y(n1150) );
  NAND2X1 U1854 ( .A(\mem<0><4> ), .B(n45), .Y(n1833) );
  OAI21X1 U1855 ( .A(n1269), .B(n1283), .C(n1833), .Y(n1151) );
  NAND2X1 U1856 ( .A(\mem<0><5> ), .B(n45), .Y(n1834) );
  OAI21X1 U1857 ( .A(n1269), .B(n1285), .C(n1834), .Y(n1152) );
  NAND2X1 U1858 ( .A(\mem<0><6> ), .B(n45), .Y(n1835) );
  OAI21X1 U1859 ( .A(n1269), .B(n1287), .C(n1835), .Y(n1153) );
  NAND2X1 U1860 ( .A(\mem<0><7> ), .B(n45), .Y(n1836) );
  OAI21X1 U1861 ( .A(n1269), .B(n1289), .C(n1836), .Y(n1154) );
  NAND2X1 U1862 ( .A(\mem<0><8> ), .B(n45), .Y(n1837) );
  OAI21X1 U1863 ( .A(n1269), .B(n1291), .C(n1837), .Y(n1155) );
  NAND2X1 U1864 ( .A(\mem<0><9> ), .B(n45), .Y(n1838) );
  OAI21X1 U1865 ( .A(n1269), .B(n1293), .C(n1838), .Y(n1156) );
  NAND2X1 U1866 ( .A(\mem<0><10> ), .B(n45), .Y(n1839) );
  OAI21X1 U1867 ( .A(n1269), .B(n1295), .C(n1839), .Y(n1157) );
  NAND2X1 U1868 ( .A(\mem<0><11> ), .B(n45), .Y(n1840) );
  OAI21X1 U1869 ( .A(n1269), .B(n1297), .C(n1840), .Y(n1158) );
  NAND2X1 U1870 ( .A(\mem<0><12> ), .B(n45), .Y(n1841) );
  OAI21X1 U1871 ( .A(n1269), .B(n1299), .C(n1841), .Y(n1159) );
  NAND2X1 U1872 ( .A(\mem<0><13> ), .B(n45), .Y(n1842) );
  OAI21X1 U1873 ( .A(n1269), .B(n1301), .C(n1842), .Y(n1160) );
  NAND2X1 U1874 ( .A(\mem<0><14> ), .B(n45), .Y(n1843) );
  OAI21X1 U1875 ( .A(n1269), .B(n1303), .C(n1843), .Y(n1161) );
  NAND2X1 U1876 ( .A(\mem<0><15> ), .B(n45), .Y(n1844) );
  OAI21X1 U1877 ( .A(n1269), .B(n1305), .C(n1844), .Y(n1162) );
endmodule


module memc_Size16_2 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n1833), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n1834), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n1835), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n1836), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n1837), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n1838), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n1839), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n1840), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n1841), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1842), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1843), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1844), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1845), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1846), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1847), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1848), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n1849), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n1850), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n1851), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n1852), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n1853), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n1854), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n1855), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n1856), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1857), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1858), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1859), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1860), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1861), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1862), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1863), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1864), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n1865), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n1866), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n1867), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n1868), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n1869), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n1870), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n1871), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n1872), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1873), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1874), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1875), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1876), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1877), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1878), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1879), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1880), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n1881), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n1882), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n1883), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n1884), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n1885), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n1886), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n1887), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n1888), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1889), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1890), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1891), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1892), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1893), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1894), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1895), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1896), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n1897), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n1898), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n1899), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n1900), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n1901), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n1902), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n1903), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n1904), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1905), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1906), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1907), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1908), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1909), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1910), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1911), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1912), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n1913), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n1914), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n1915), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n1916), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n1917), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n1918), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n1919), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n1920), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1921), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1922), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1923), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1924), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1925), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1926), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1927), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1928), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n1929), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n1930), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n1931), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n1932), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n1933), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n1934), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n1935), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n1936), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1937), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1938), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1939), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1940), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1941), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1942), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1943), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1944), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n1945), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n1946), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n1947), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n1948), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n1949), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n1950), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n1951), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n1952), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1953), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1954), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1955), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1956), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1957), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1958), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1959), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1960), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n1961), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n1962), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n1963), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n1964), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n1965), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n1966), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n1967), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n1968), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1969), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1970), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1971), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1972), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1973), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1974), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1975), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1976), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n1977), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n1978), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n1979), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n1980), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n1981), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n1982), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n1983), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n1984), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n1985), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n1986), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n1987), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n1988), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n1989), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n1990), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n1991), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n1992), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n1993), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n1994), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n1995), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n1996), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n1997), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n1998), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n1999), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n2000), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n2001), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n2002), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n2003), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n2004), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n2005), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n2006), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n2007), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n2008), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n2009), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n2010), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n2011), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n2012), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n2013), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n2014), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n2015), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n2016), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n2017), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n2018), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n2019), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n2020), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n2021), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n2022), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n2023), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n2024), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n2025), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n2026), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n2027), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n2028), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n2029), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n2030), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n2031), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n2032), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2033), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2034), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2035), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2036), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2037), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2038), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2039), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2040), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n2041), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n2042), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n2043), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n2044), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n2045), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n2046), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n2047), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n2048), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2049), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2050), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2051), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2052), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2053), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2054), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2055), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2056), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n2057), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n2058), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n2059), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n2060), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n2061), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n2062), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n2063), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n2064), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2065), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2066), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2067), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2068), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2069), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2070), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2071), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2072), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n2073), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n2074), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n2075), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n2076), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n2077), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n2078), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n2079), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n2080), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2081), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2082), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2083), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2084), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2085), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2086), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2087), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2088), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n2089), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n2090), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n2091), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n2092), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n2093), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n2094), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n2095), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n2096), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2097), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2098), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2099), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2100), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2101), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2102), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2103), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2104), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n2105), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n2106), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n2107), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n2108), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n2109), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n2110), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n2111), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n2112), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2113), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2114), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2115), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2116), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2117), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2118), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2119), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2120), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n2121), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n2122), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n2123), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n2124), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n2125), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n2126), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n2127), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n2128), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2129), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2130), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2131), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2132), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2133), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2134), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2135), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2136), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n2137), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n2138), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n2139), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n2140), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n2141), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n2142), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n2143), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n2144), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2145), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2146), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2147), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2148), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2149), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2150), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2151), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2152), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n2153), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n2154), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n2155), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n2156), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n2157), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n2158), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n2159), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n2160), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2161), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2162), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2163), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2164), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2165), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2166), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2167), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2168), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n2169), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n2170), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n2171), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n2172), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n2173), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n2174), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n2175), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n2176), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2177), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2178), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2179), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2180), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2181), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2182), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2183), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2184), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n2185), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n2186), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n2187), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n2188), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n2189), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n2190), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n2191), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n2192), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2193), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2194), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2195), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2196), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2197), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2198), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2199), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2200), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n2201), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n2202), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n2203), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n2204), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n2205), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n2206), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n2207), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n2208), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2209), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2210), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2211), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2212), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2213), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2214), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2215), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2216), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n2217), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n2218), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n2219), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n2220), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n2221), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n2222), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n2223), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n2224), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2225), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2226), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2227), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2228), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2229), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2230), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2231), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2232), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n2233), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n2234), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n2235), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n2236), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n2237), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n2238), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n2239), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n2240), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2241), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2242), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2243), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2244), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2245), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2246), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2247), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2248), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n2249), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n2250), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n2251), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n2252), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n2253), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n2254), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n2255), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n2256), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2257), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2258), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2259), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2260), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2261), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2262), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2263), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2264), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n2265), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n2266), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n2267), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n2268), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n2269), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n2270), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n2271), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n2272), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2273), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2274), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2275), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2276), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2277), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2278), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2279), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2280), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n2281), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n2282), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n2283), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n2284), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n2285), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n2286), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n2287), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n2288), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2289), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2290), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2291), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2292), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2293), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2294), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2295), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2296), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n2297), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n2298), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n2299), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n2300), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n2301), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n2302), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n2303), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n2304), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2305), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2306), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2307), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2308), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2309), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2310), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2311), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2312), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n2313), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n2314), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n2315), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n2316), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n2317), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n2318), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n2319), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n2320), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2321), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2322), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2323), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2324), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2325), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2326), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2327), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2328), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n2329), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n2330), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n2331), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n2332), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n2333), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n2334), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n2335), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n2336), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2337), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2338), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2339), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2340), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2341), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2342), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2343), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2344), .CLK(clk), .Q(\mem<31><0> ) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n2345) );
  INVX1 U2 ( .A(n1211), .Y(n1192) );
  INVX2 U3 ( .A(N10), .Y(n1295) );
  INVX2 U4 ( .A(n1192), .Y(n1198) );
  INVX2 U5 ( .A(n1192), .Y(n1200) );
  INVX2 U6 ( .A(n1192), .Y(n1199) );
  INVX2 U7 ( .A(n1192), .Y(n1207) );
  INVX2 U8 ( .A(n1192), .Y(n1208) );
  INVX1 U9 ( .A(n1295), .Y(n1202) );
  INVX1 U10 ( .A(n1295), .Y(n1204) );
  INVX1 U11 ( .A(n1295), .Y(n1201) );
  INVX1 U12 ( .A(n1295), .Y(n1205) );
  INVX1 U13 ( .A(n1193), .Y(n1203) );
  INVX1 U14 ( .A(n1295), .Y(n1206) );
  INVX1 U15 ( .A(n1295), .Y(n1209) );
  INVX4 U16 ( .A(n51), .Y(n140) );
  INVX4 U17 ( .A(n50), .Y(n137) );
  AND2X2 U18 ( .A(n1295), .B(n60), .Y(n71) );
  INVX1 U19 ( .A(n644), .Y(N30) );
  INVX2 U20 ( .A(n1193), .Y(n1194) );
  INVX1 U21 ( .A(n1191), .Y(n1180) );
  INVX2 U22 ( .A(n1193), .Y(n1195) );
  INVX1 U23 ( .A(n1191), .Y(n1181) );
  INVX1 U24 ( .A(n1192), .Y(n1197) );
  INVX1 U25 ( .A(n1193), .Y(n1196) );
  INVX1 U26 ( .A(n1191), .Y(n1182) );
  INVX1 U27 ( .A(n1179), .Y(n1183) );
  INVX1 U28 ( .A(n1179), .Y(n1184) );
  INVX1 U29 ( .A(n1179), .Y(n1185) );
  INVX1 U30 ( .A(n1178), .Y(n1186) );
  INVX1 U31 ( .A(n1178), .Y(n1187) );
  INVX1 U32 ( .A(n1178), .Y(n1188) );
  INVX1 U33 ( .A(n1179), .Y(n1189) );
  INVX1 U34 ( .A(n1178), .Y(n1190) );
  INVX1 U35 ( .A(n1301), .Y(n1173) );
  INVX1 U36 ( .A(n1301), .Y(n1172) );
  INVX1 U37 ( .A(n1301), .Y(n1171) );
  INVX1 U38 ( .A(n642), .Y(N32) );
  INVX1 U39 ( .A(n643), .Y(N31) );
  INVX1 U40 ( .A(n645), .Y(N29) );
  INVX1 U41 ( .A(n646), .Y(N28) );
  INVX1 U42 ( .A(n647), .Y(N27) );
  INVX1 U43 ( .A(n648), .Y(N26) );
  INVX1 U44 ( .A(n649), .Y(N25) );
  INVX1 U45 ( .A(n650), .Y(N24) );
  INVX1 U46 ( .A(n1163), .Y(N23) );
  INVX1 U47 ( .A(n1164), .Y(N22) );
  INVX1 U48 ( .A(n1165), .Y(N21) );
  INVX1 U49 ( .A(n1166), .Y(N20) );
  INVX1 U50 ( .A(n1167), .Y(N19) );
  INVX1 U51 ( .A(n1168), .Y(N18) );
  INVX1 U52 ( .A(n1169), .Y(N17) );
  INVX1 U53 ( .A(n1299), .Y(n1176) );
  INVX1 U54 ( .A(n1299), .Y(n1177) );
  INVX1 U55 ( .A(n1296), .Y(n1191) );
  INVX1 U56 ( .A(n1299), .Y(n1175) );
  INVX1 U57 ( .A(n1299), .Y(n1174) );
  INVX1 U58 ( .A(n1295), .Y(n1211) );
  INVX1 U59 ( .A(N14), .Y(n1303) );
  INVX1 U60 ( .A(n1211), .Y(n1193) );
  INVX2 U61 ( .A(n1192), .Y(n1210) );
  INVX1 U62 ( .A(n1296), .Y(n1178) );
  INVX1 U63 ( .A(n1296), .Y(n1179) );
  INVX1 U64 ( .A(n1303), .Y(n1170) );
  INVX1 U65 ( .A(rst), .Y(n1294) );
  INVX1 U66 ( .A(n89), .Y(n1226) );
  INVX1 U67 ( .A(n90), .Y(n1243) );
  INVX1 U68 ( .A(n91), .Y(n1260) );
  INVX1 U69 ( .A(n92), .Y(n1263) );
  INVX2 U70 ( .A(n1304), .Y(n1305) );
  INVX1 U71 ( .A(N13), .Y(n1301) );
  INVX2 U72 ( .A(n1304), .Y(n1) );
  AND2X2 U73 ( .A(n1266), .B(n93), .Y(n2) );
  INVX1 U74 ( .A(n2), .Y(n3) );
  AND2X2 U75 ( .A(n1268), .B(n95), .Y(n4) );
  INVX1 U76 ( .A(n4), .Y(n5) );
  AND2X2 U77 ( .A(n1266), .B(n97), .Y(n6) );
  INVX1 U78 ( .A(n6), .Y(n7) );
  AND2X2 U79 ( .A(n1268), .B(n99), .Y(n8) );
  INVX1 U80 ( .A(n8), .Y(n9) );
  AND2X2 U81 ( .A(n1266), .B(n101), .Y(n10) );
  INVX1 U82 ( .A(n10), .Y(n11) );
  AND2X2 U83 ( .A(n1268), .B(n103), .Y(n12) );
  INVX1 U84 ( .A(n12), .Y(n13) );
  AND2X2 U85 ( .A(n1267), .B(n105), .Y(n14) );
  INVX1 U86 ( .A(n14), .Y(n15) );
  AND2X2 U87 ( .A(n1268), .B(n89), .Y(n16) );
  INVX1 U88 ( .A(n16), .Y(n17) );
  AND2X2 U89 ( .A(n1266), .B(n107), .Y(n18) );
  INVX1 U90 ( .A(n18), .Y(n19) );
  AND2X2 U91 ( .A(n1268), .B(n109), .Y(n20) );
  INVX1 U92 ( .A(n20), .Y(n21) );
  AND2X2 U93 ( .A(n1267), .B(n111), .Y(n22) );
  INVX1 U94 ( .A(n22), .Y(n23) );
  AND2X2 U95 ( .A(n1266), .B(n113), .Y(n24) );
  INVX1 U96 ( .A(n24), .Y(n25) );
  AND2X2 U97 ( .A(n1266), .B(n115), .Y(n26) );
  INVX1 U98 ( .A(n26), .Y(n27) );
  AND2X2 U99 ( .A(n1266), .B(n117), .Y(n28) );
  INVX1 U100 ( .A(n28), .Y(n29) );
  AND2X2 U101 ( .A(n1266), .B(n119), .Y(n30) );
  INVX1 U102 ( .A(n30), .Y(n31) );
  AND2X2 U103 ( .A(n1266), .B(n90), .Y(n32) );
  INVX1 U104 ( .A(n32), .Y(n33) );
  AND2X2 U105 ( .A(n1266), .B(n121), .Y(n34) );
  INVX1 U106 ( .A(n34), .Y(n35) );
  AND2X2 U107 ( .A(n1266), .B(n123), .Y(n36) );
  INVX1 U108 ( .A(n36), .Y(n37) );
  AND2X2 U109 ( .A(n1266), .B(n125), .Y(n38) );
  INVX1 U110 ( .A(n38), .Y(n39) );
  AND2X2 U111 ( .A(n1266), .B(n127), .Y(n40) );
  INVX1 U112 ( .A(n40), .Y(n41) );
  AND2X2 U113 ( .A(n1266), .B(n129), .Y(n42) );
  INVX1 U114 ( .A(n42), .Y(n43) );
  AND2X2 U115 ( .A(n1266), .B(n131), .Y(n44) );
  INVX1 U116 ( .A(n44), .Y(n45) );
  AND2X2 U117 ( .A(n1266), .B(n133), .Y(n46) );
  INVX1 U118 ( .A(n46), .Y(n47) );
  AND2X2 U119 ( .A(n1267), .B(n91), .Y(n48) );
  INVX1 U120 ( .A(n48), .Y(n49) );
  AND2X2 U121 ( .A(n1267), .B(n135), .Y(n50) );
  AND2X2 U122 ( .A(n1267), .B(n138), .Y(n51) );
  AND2X2 U123 ( .A(n1267), .B(n141), .Y(n52) );
  AND2X2 U124 ( .A(n1267), .B(n145), .Y(n53) );
  AND2X2 U125 ( .A(n1267), .B(n149), .Y(n54) );
  AND2X2 U126 ( .A(n1267), .B(n153), .Y(n55) );
  AND2X2 U127 ( .A(n1267), .B(n157), .Y(n56) );
  AND2X2 U128 ( .A(n1266), .B(n92), .Y(n57) );
  INVX1 U129 ( .A(n57), .Y(n58) );
  BUFX2 U130 ( .A(n3), .Y(n1212) );
  BUFX2 U131 ( .A(n3), .Y(n1213) );
  BUFX2 U132 ( .A(n5), .Y(n1214) );
  BUFX2 U133 ( .A(n5), .Y(n1215) );
  BUFX2 U134 ( .A(n7), .Y(n1216) );
  BUFX2 U135 ( .A(n7), .Y(n1217) );
  BUFX2 U136 ( .A(n9), .Y(n1218) );
  BUFX2 U137 ( .A(n9), .Y(n1219) );
  BUFX2 U138 ( .A(n11), .Y(n1220) );
  BUFX2 U139 ( .A(n11), .Y(n1221) );
  BUFX2 U140 ( .A(n13), .Y(n1222) );
  BUFX2 U141 ( .A(n13), .Y(n1223) );
  BUFX2 U142 ( .A(n15), .Y(n1224) );
  BUFX2 U143 ( .A(n15), .Y(n1225) );
  BUFX2 U144 ( .A(n17), .Y(n1227) );
  BUFX2 U145 ( .A(n17), .Y(n1228) );
  BUFX2 U146 ( .A(n19), .Y(n1229) );
  BUFX2 U147 ( .A(n19), .Y(n1230) );
  BUFX2 U148 ( .A(n21), .Y(n1231) );
  BUFX2 U149 ( .A(n21), .Y(n1232) );
  BUFX2 U150 ( .A(n23), .Y(n1233) );
  BUFX2 U151 ( .A(n23), .Y(n1234) );
  BUFX2 U152 ( .A(n25), .Y(n1235) );
  BUFX2 U153 ( .A(n25), .Y(n1236) );
  BUFX2 U154 ( .A(n27), .Y(n1237) );
  BUFX2 U155 ( .A(n27), .Y(n1238) );
  BUFX2 U156 ( .A(n29), .Y(n1239) );
  BUFX2 U157 ( .A(n29), .Y(n1240) );
  BUFX2 U158 ( .A(n31), .Y(n1241) );
  BUFX2 U159 ( .A(n31), .Y(n1242) );
  BUFX2 U160 ( .A(n33), .Y(n1244) );
  BUFX2 U161 ( .A(n33), .Y(n1245) );
  BUFX2 U162 ( .A(n35), .Y(n1246) );
  BUFX2 U163 ( .A(n35), .Y(n1247) );
  BUFX2 U164 ( .A(n37), .Y(n1248) );
  BUFX2 U165 ( .A(n37), .Y(n1249) );
  BUFX2 U166 ( .A(n39), .Y(n1250) );
  BUFX2 U167 ( .A(n39), .Y(n1251) );
  BUFX2 U168 ( .A(n41), .Y(n1252) );
  BUFX2 U169 ( .A(n41), .Y(n1253) );
  BUFX2 U170 ( .A(n43), .Y(n1254) );
  BUFX2 U171 ( .A(n43), .Y(n1255) );
  BUFX2 U172 ( .A(n45), .Y(n1256) );
  BUFX2 U173 ( .A(n45), .Y(n1257) );
  BUFX2 U174 ( .A(n47), .Y(n1258) );
  BUFX2 U175 ( .A(n47), .Y(n1259) );
  BUFX2 U176 ( .A(n49), .Y(n1261) );
  BUFX2 U177 ( .A(n49), .Y(n1262) );
  BUFX2 U178 ( .A(n58), .Y(n1264) );
  BUFX2 U179 ( .A(n58), .Y(n1265) );
  AND2X2 U180 ( .A(write), .B(n1294), .Y(n59) );
  INVX1 U181 ( .A(n1297), .Y(n1296) );
  INVX1 U182 ( .A(n1301), .Y(n1300) );
  AND2X1 U183 ( .A(n1298), .B(n1296), .Y(n60) );
  INVX1 U184 ( .A(n1299), .Y(n1298) );
  AND2X1 U185 ( .A(n2345), .B(n1302), .Y(n61) );
  INVX1 U186 ( .A(n1303), .Y(n1302) );
  BUFX2 U187 ( .A(n1338), .Y(n62) );
  INVX1 U188 ( .A(n62), .Y(n1730) );
  BUFX2 U189 ( .A(n1355), .Y(n63) );
  INVX1 U190 ( .A(n63), .Y(n1747) );
  BUFX2 U191 ( .A(n1372), .Y(n64) );
  INVX1 U192 ( .A(n64), .Y(n1764) );
  BUFX2 U193 ( .A(n1389), .Y(n65) );
  INVX1 U194 ( .A(n65), .Y(n1781) );
  BUFX2 U195 ( .A(n1406), .Y(n66) );
  INVX1 U196 ( .A(n66), .Y(n1798) );
  BUFX2 U197 ( .A(n1567), .Y(n67) );
  INVX1 U198 ( .A(n67), .Y(n1680) );
  BUFX2 U199 ( .A(n1697), .Y(n68) );
  INVX1 U200 ( .A(n68), .Y(n1815) );
  AND2X1 U201 ( .A(N10), .B(n60), .Y(n69) );
  AND2X1 U202 ( .A(n1300), .B(n61), .Y(n70) );
  AND2X1 U203 ( .A(n1301), .B(n61), .Y(n72) );
  AND2X2 U204 ( .A(\data_in<0> ), .B(n1268), .Y(n73) );
  AND2X2 U205 ( .A(\data_in<1> ), .B(n1268), .Y(n74) );
  AND2X2 U206 ( .A(\data_in<2> ), .B(n1268), .Y(n75) );
  AND2X2 U207 ( .A(\data_in<3> ), .B(n1268), .Y(n76) );
  AND2X2 U208 ( .A(\data_in<4> ), .B(n1268), .Y(n77) );
  AND2X2 U209 ( .A(\data_in<5> ), .B(n1268), .Y(n78) );
  AND2X2 U210 ( .A(\data_in<6> ), .B(n1268), .Y(n79) );
  AND2X2 U211 ( .A(\data_in<7> ), .B(n1268), .Y(n80) );
  AND2X2 U212 ( .A(\data_in<8> ), .B(n1268), .Y(n81) );
  AND2X2 U213 ( .A(\data_in<9> ), .B(n1268), .Y(n82) );
  AND2X2 U214 ( .A(\data_in<10> ), .B(n1268), .Y(n83) );
  AND2X2 U215 ( .A(\data_in<11> ), .B(n1267), .Y(n84) );
  AND2X2 U216 ( .A(\data_in<12> ), .B(n1267), .Y(n85) );
  AND2X2 U217 ( .A(\data_in<13> ), .B(n1267), .Y(n86) );
  AND2X2 U218 ( .A(\data_in<14> ), .B(n1267), .Y(n87) );
  AND2X2 U219 ( .A(\data_in<15> ), .B(n1267), .Y(n88) );
  AND2X1 U220 ( .A(n70), .B(n1816), .Y(n89) );
  AND2X1 U221 ( .A(n1816), .B(n72), .Y(n90) );
  AND2X1 U222 ( .A(n1816), .B(n1680), .Y(n91) );
  AND2X1 U223 ( .A(n1816), .B(n1815), .Y(n92) );
  AND2X1 U224 ( .A(n69), .B(n70), .Y(n93) );
  INVX1 U225 ( .A(n93), .Y(n94) );
  AND2X1 U226 ( .A(n70), .B(n71), .Y(n95) );
  INVX1 U227 ( .A(n95), .Y(n96) );
  AND2X1 U228 ( .A(n70), .B(n1730), .Y(n97) );
  INVX1 U229 ( .A(n97), .Y(n98) );
  AND2X1 U230 ( .A(n70), .B(n1747), .Y(n99) );
  INVX1 U231 ( .A(n99), .Y(n100) );
  AND2X1 U232 ( .A(n70), .B(n1764), .Y(n101) );
  INVX1 U233 ( .A(n101), .Y(n102) );
  AND2X1 U234 ( .A(n70), .B(n1781), .Y(n103) );
  INVX1 U235 ( .A(n103), .Y(n104) );
  AND2X1 U236 ( .A(n70), .B(n1798), .Y(n105) );
  INVX1 U237 ( .A(n105), .Y(n106) );
  AND2X1 U238 ( .A(n69), .B(n72), .Y(n107) );
  INVX1 U239 ( .A(n107), .Y(n108) );
  AND2X1 U240 ( .A(n71), .B(n72), .Y(n109) );
  INVX1 U241 ( .A(n109), .Y(n110) );
  AND2X1 U242 ( .A(n1730), .B(n72), .Y(n111) );
  INVX1 U243 ( .A(n111), .Y(n112) );
  AND2X1 U244 ( .A(n1747), .B(n72), .Y(n113) );
  INVX1 U245 ( .A(n113), .Y(n114) );
  AND2X1 U246 ( .A(n1764), .B(n72), .Y(n115) );
  INVX1 U247 ( .A(n115), .Y(n116) );
  AND2X1 U248 ( .A(n1781), .B(n72), .Y(n117) );
  INVX1 U249 ( .A(n117), .Y(n118) );
  AND2X1 U250 ( .A(n1798), .B(n72), .Y(n119) );
  INVX1 U251 ( .A(n119), .Y(n120) );
  AND2X1 U252 ( .A(n69), .B(n1680), .Y(n121) );
  INVX1 U253 ( .A(n121), .Y(n122) );
  AND2X1 U254 ( .A(n71), .B(n1680), .Y(n123) );
  INVX1 U255 ( .A(n123), .Y(n124) );
  AND2X1 U256 ( .A(n1730), .B(n1680), .Y(n125) );
  INVX1 U257 ( .A(n125), .Y(n126) );
  AND2X1 U258 ( .A(n1747), .B(n1680), .Y(n127) );
  INVX1 U259 ( .A(n127), .Y(n128) );
  AND2X1 U260 ( .A(n1764), .B(n1680), .Y(n129) );
  INVX1 U261 ( .A(n129), .Y(n130) );
  AND2X1 U262 ( .A(n1781), .B(n1680), .Y(n131) );
  INVX1 U263 ( .A(n131), .Y(n132) );
  AND2X1 U264 ( .A(n1798), .B(n1680), .Y(n133) );
  INVX1 U265 ( .A(n133), .Y(n134) );
  AND2X1 U266 ( .A(n69), .B(n1815), .Y(n135) );
  INVX1 U267 ( .A(n135), .Y(n136) );
  AND2X1 U268 ( .A(n71), .B(n1815), .Y(n138) );
  INVX1 U269 ( .A(n138), .Y(n139) );
  AND2X1 U270 ( .A(n1730), .B(n1815), .Y(n141) );
  INVX1 U271 ( .A(n141), .Y(n142) );
  INVX1 U272 ( .A(n52), .Y(n143) );
  INVX1 U273 ( .A(n52), .Y(n144) );
  AND2X1 U274 ( .A(n1747), .B(n1815), .Y(n145) );
  INVX1 U275 ( .A(n145), .Y(n146) );
  INVX1 U276 ( .A(n53), .Y(n147) );
  INVX1 U277 ( .A(n53), .Y(n148) );
  AND2X1 U278 ( .A(n1764), .B(n1815), .Y(n149) );
  INVX1 U279 ( .A(n149), .Y(n150) );
  INVX1 U280 ( .A(n54), .Y(n151) );
  INVX1 U281 ( .A(n54), .Y(n152) );
  AND2X1 U282 ( .A(n1781), .B(n1815), .Y(n153) );
  INVX1 U283 ( .A(n153), .Y(n154) );
  INVX1 U284 ( .A(n55), .Y(n155) );
  INVX1 U285 ( .A(n55), .Y(n156) );
  AND2X1 U286 ( .A(n1798), .B(n1815), .Y(n157) );
  INVX1 U287 ( .A(n157), .Y(n158) );
  INVX1 U288 ( .A(n56), .Y(n159) );
  INVX1 U289 ( .A(n56), .Y(n160) );
  MUX2X1 U290 ( .B(n162), .A(n163), .S(n1180), .Y(n161) );
  MUX2X1 U291 ( .B(n165), .A(n166), .S(n1180), .Y(n164) );
  MUX2X1 U292 ( .B(n168), .A(n169), .S(n1180), .Y(n167) );
  MUX2X1 U293 ( .B(n171), .A(n172), .S(n1180), .Y(n170) );
  MUX2X1 U294 ( .B(n174), .A(n175), .S(n1173), .Y(n173) );
  MUX2X1 U295 ( .B(n177), .A(n178), .S(n1180), .Y(n176) );
  MUX2X1 U296 ( .B(n180), .A(n181), .S(n1180), .Y(n179) );
  MUX2X1 U297 ( .B(n183), .A(n184), .S(n1180), .Y(n182) );
  MUX2X1 U298 ( .B(n186), .A(n187), .S(n1180), .Y(n185) );
  MUX2X1 U299 ( .B(n189), .A(n190), .S(n1173), .Y(n188) );
  MUX2X1 U300 ( .B(n192), .A(n193), .S(n1181), .Y(n191) );
  MUX2X1 U301 ( .B(n195), .A(n196), .S(n1181), .Y(n194) );
  MUX2X1 U302 ( .B(n198), .A(n199), .S(n1181), .Y(n197) );
  MUX2X1 U303 ( .B(n201), .A(n202), .S(n1181), .Y(n200) );
  MUX2X1 U304 ( .B(n204), .A(n205), .S(n1173), .Y(n203) );
  MUX2X1 U305 ( .B(n207), .A(n208), .S(n1181), .Y(n206) );
  MUX2X1 U306 ( .B(n210), .A(n211), .S(n1181), .Y(n209) );
  MUX2X1 U307 ( .B(n213), .A(n215), .S(n1181), .Y(n212) );
  MUX2X1 U308 ( .B(n217), .A(n218), .S(n1181), .Y(n216) );
  MUX2X1 U309 ( .B(n220), .A(n221), .S(n1173), .Y(n219) );
  MUX2X1 U310 ( .B(n223), .A(n224), .S(n1181), .Y(n222) );
  MUX2X1 U311 ( .B(n226), .A(n227), .S(n1181), .Y(n225) );
  MUX2X1 U312 ( .B(n229), .A(n230), .S(n1181), .Y(n228) );
  MUX2X1 U313 ( .B(n232), .A(n233), .S(n1181), .Y(n231) );
  MUX2X1 U314 ( .B(n235), .A(n236), .S(n1173), .Y(n234) );
  MUX2X1 U315 ( .B(n238), .A(n239), .S(n1182), .Y(n237) );
  MUX2X1 U316 ( .B(n241), .A(n242), .S(n1182), .Y(n240) );
  MUX2X1 U317 ( .B(n244), .A(n245), .S(n1182), .Y(n243) );
  MUX2X1 U318 ( .B(n247), .A(n248), .S(n1182), .Y(n246) );
  MUX2X1 U319 ( .B(n250), .A(n251), .S(n1173), .Y(n249) );
  MUX2X1 U320 ( .B(n253), .A(n254), .S(n1182), .Y(n252) );
  MUX2X1 U321 ( .B(n256), .A(n257), .S(n1182), .Y(n255) );
  MUX2X1 U322 ( .B(n259), .A(n260), .S(n1182), .Y(n258) );
  MUX2X1 U323 ( .B(n262), .A(n263), .S(n1182), .Y(n261) );
  MUX2X1 U324 ( .B(n265), .A(n266), .S(n1173), .Y(n264) );
  MUX2X1 U325 ( .B(n268), .A(n269), .S(n1182), .Y(n267) );
  MUX2X1 U326 ( .B(n271), .A(n272), .S(n1182), .Y(n270) );
  MUX2X1 U327 ( .B(n274), .A(n275), .S(n1182), .Y(n273) );
  MUX2X1 U328 ( .B(n277), .A(n278), .S(n1182), .Y(n276) );
  MUX2X1 U329 ( .B(n280), .A(n281), .S(n1173), .Y(n279) );
  MUX2X1 U330 ( .B(n283), .A(n284), .S(n1183), .Y(n282) );
  MUX2X1 U331 ( .B(n286), .A(n287), .S(n1183), .Y(n285) );
  MUX2X1 U332 ( .B(n289), .A(n290), .S(n1183), .Y(n288) );
  MUX2X1 U333 ( .B(n292), .A(n293), .S(n1183), .Y(n291) );
  MUX2X1 U334 ( .B(n295), .A(n296), .S(n1173), .Y(n294) );
  MUX2X1 U335 ( .B(n298), .A(n299), .S(n1183), .Y(n297) );
  MUX2X1 U336 ( .B(n301), .A(n302), .S(n1183), .Y(n300) );
  MUX2X1 U337 ( .B(n304), .A(n305), .S(n1183), .Y(n303) );
  MUX2X1 U338 ( .B(n307), .A(n308), .S(n1183), .Y(n306) );
  MUX2X1 U339 ( .B(n310), .A(n311), .S(n1173), .Y(n309) );
  MUX2X1 U340 ( .B(n313), .A(n314), .S(n1183), .Y(n312) );
  MUX2X1 U341 ( .B(n316), .A(n317), .S(n1183), .Y(n315) );
  MUX2X1 U342 ( .B(n319), .A(n320), .S(n1183), .Y(n318) );
  MUX2X1 U343 ( .B(n322), .A(n323), .S(n1183), .Y(n321) );
  MUX2X1 U344 ( .B(n325), .A(n326), .S(n1173), .Y(n324) );
  MUX2X1 U345 ( .B(n328), .A(n329), .S(n1184), .Y(n327) );
  MUX2X1 U346 ( .B(n331), .A(n332), .S(n1184), .Y(n330) );
  MUX2X1 U347 ( .B(n334), .A(n335), .S(n1184), .Y(n333) );
  MUX2X1 U348 ( .B(n337), .A(n338), .S(n1184), .Y(n336) );
  MUX2X1 U349 ( .B(n340), .A(n341), .S(n1173), .Y(n339) );
  MUX2X1 U350 ( .B(n343), .A(n344), .S(n1184), .Y(n342) );
  MUX2X1 U351 ( .B(n346), .A(n347), .S(n1184), .Y(n345) );
  MUX2X1 U352 ( .B(n349), .A(n350), .S(n1184), .Y(n348) );
  MUX2X1 U353 ( .B(n352), .A(n353), .S(n1184), .Y(n351) );
  MUX2X1 U354 ( .B(n355), .A(n356), .S(n1172), .Y(n354) );
  MUX2X1 U355 ( .B(n358), .A(n359), .S(n1184), .Y(n357) );
  MUX2X1 U356 ( .B(n361), .A(n362), .S(n1184), .Y(n360) );
  MUX2X1 U357 ( .B(n364), .A(n365), .S(n1184), .Y(n363) );
  MUX2X1 U358 ( .B(n367), .A(n368), .S(n1184), .Y(n366) );
  MUX2X1 U359 ( .B(n370), .A(n371), .S(n1172), .Y(n369) );
  MUX2X1 U360 ( .B(n373), .A(n374), .S(n1185), .Y(n372) );
  MUX2X1 U361 ( .B(n376), .A(n377), .S(n1185), .Y(n375) );
  MUX2X1 U362 ( .B(n379), .A(n380), .S(n1185), .Y(n378) );
  MUX2X1 U363 ( .B(n382), .A(n383), .S(n1185), .Y(n381) );
  MUX2X1 U364 ( .B(n385), .A(n386), .S(n1172), .Y(n384) );
  MUX2X1 U365 ( .B(n388), .A(n389), .S(n1185), .Y(n387) );
  MUX2X1 U366 ( .B(n391), .A(n392), .S(n1185), .Y(n390) );
  MUX2X1 U367 ( .B(n394), .A(n395), .S(n1185), .Y(n393) );
  MUX2X1 U368 ( .B(n397), .A(n398), .S(n1185), .Y(n396) );
  MUX2X1 U369 ( .B(n400), .A(n401), .S(n1172), .Y(n399) );
  MUX2X1 U370 ( .B(n403), .A(n404), .S(n1185), .Y(n402) );
  MUX2X1 U371 ( .B(n406), .A(n407), .S(n1185), .Y(n405) );
  MUX2X1 U372 ( .B(n409), .A(n410), .S(n1185), .Y(n408) );
  MUX2X1 U373 ( .B(n412), .A(n413), .S(n1185), .Y(n411) );
  MUX2X1 U374 ( .B(n415), .A(n416), .S(n1172), .Y(n414) );
  MUX2X1 U375 ( .B(n418), .A(n419), .S(n1186), .Y(n417) );
  MUX2X1 U376 ( .B(n421), .A(n422), .S(n1186), .Y(n420) );
  MUX2X1 U377 ( .B(n424), .A(n425), .S(n1186), .Y(n423) );
  MUX2X1 U378 ( .B(n427), .A(n428), .S(n1186), .Y(n426) );
  MUX2X1 U379 ( .B(n430), .A(n431), .S(n1172), .Y(n429) );
  MUX2X1 U380 ( .B(n433), .A(n434), .S(n1186), .Y(n432) );
  MUX2X1 U381 ( .B(n436), .A(n437), .S(n1186), .Y(n435) );
  MUX2X1 U382 ( .B(n439), .A(n440), .S(n1186), .Y(n438) );
  MUX2X1 U383 ( .B(n442), .A(n443), .S(n1186), .Y(n441) );
  MUX2X1 U384 ( .B(n445), .A(n446), .S(n1172), .Y(n444) );
  MUX2X1 U385 ( .B(n448), .A(n449), .S(n1186), .Y(n447) );
  MUX2X1 U386 ( .B(n451), .A(n452), .S(n1186), .Y(n450) );
  MUX2X1 U387 ( .B(n454), .A(n455), .S(n1186), .Y(n453) );
  MUX2X1 U388 ( .B(n457), .A(n458), .S(n1186), .Y(n456) );
  MUX2X1 U389 ( .B(n460), .A(n461), .S(n1172), .Y(n459) );
  MUX2X1 U390 ( .B(n463), .A(n464), .S(n1187), .Y(n462) );
  MUX2X1 U391 ( .B(n466), .A(n467), .S(n1187), .Y(n465) );
  MUX2X1 U392 ( .B(n469), .A(n470), .S(n1187), .Y(n468) );
  MUX2X1 U393 ( .B(n472), .A(n473), .S(n1187), .Y(n471) );
  MUX2X1 U394 ( .B(n475), .A(n476), .S(n1172), .Y(n474) );
  MUX2X1 U395 ( .B(n478), .A(n479), .S(n1187), .Y(n477) );
  MUX2X1 U396 ( .B(n481), .A(n482), .S(n1187), .Y(n480) );
  MUX2X1 U397 ( .B(n484), .A(n485), .S(n1187), .Y(n483) );
  MUX2X1 U398 ( .B(n487), .A(n488), .S(n1187), .Y(n486) );
  MUX2X1 U399 ( .B(n490), .A(n491), .S(n1172), .Y(n489) );
  MUX2X1 U400 ( .B(n493), .A(n494), .S(n1187), .Y(n492) );
  MUX2X1 U401 ( .B(n496), .A(n497), .S(n1187), .Y(n495) );
  MUX2X1 U402 ( .B(n499), .A(n500), .S(n1187), .Y(n498) );
  MUX2X1 U403 ( .B(n502), .A(n503), .S(n1187), .Y(n501) );
  MUX2X1 U404 ( .B(n505), .A(n506), .S(n1172), .Y(n504) );
  MUX2X1 U405 ( .B(n508), .A(n509), .S(n1188), .Y(n507) );
  MUX2X1 U406 ( .B(n511), .A(n512), .S(n1188), .Y(n510) );
  MUX2X1 U407 ( .B(n514), .A(n515), .S(n1188), .Y(n513) );
  MUX2X1 U408 ( .B(n517), .A(n518), .S(n1188), .Y(n516) );
  MUX2X1 U409 ( .B(n520), .A(n521), .S(n1172), .Y(n519) );
  MUX2X1 U410 ( .B(n523), .A(n524), .S(n1188), .Y(n522) );
  MUX2X1 U411 ( .B(n526), .A(n527), .S(n1188), .Y(n525) );
  MUX2X1 U412 ( .B(n529), .A(n530), .S(n1188), .Y(n528) );
  MUX2X1 U413 ( .B(n532), .A(n533), .S(n1188), .Y(n531) );
  MUX2X1 U414 ( .B(n535), .A(n536), .S(n1171), .Y(n534) );
  MUX2X1 U415 ( .B(n538), .A(n539), .S(n1188), .Y(n537) );
  MUX2X1 U416 ( .B(n541), .A(n542), .S(n1188), .Y(n540) );
  MUX2X1 U417 ( .B(n544), .A(n545), .S(n1188), .Y(n543) );
  MUX2X1 U418 ( .B(n547), .A(n548), .S(n1188), .Y(n546) );
  MUX2X1 U419 ( .B(n550), .A(n551), .S(n1171), .Y(n549) );
  MUX2X1 U420 ( .B(n553), .A(n554), .S(n1189), .Y(n552) );
  MUX2X1 U421 ( .B(n556), .A(n557), .S(n1189), .Y(n555) );
  MUX2X1 U422 ( .B(n559), .A(n560), .S(n1189), .Y(n558) );
  MUX2X1 U423 ( .B(n562), .A(n563), .S(n1189), .Y(n561) );
  MUX2X1 U424 ( .B(n565), .A(n566), .S(n1171), .Y(n564) );
  MUX2X1 U425 ( .B(n568), .A(n569), .S(n1189), .Y(n567) );
  MUX2X1 U426 ( .B(n571), .A(n572), .S(n1189), .Y(n570) );
  MUX2X1 U427 ( .B(n574), .A(n575), .S(n1189), .Y(n573) );
  MUX2X1 U428 ( .B(n577), .A(n578), .S(n1189), .Y(n576) );
  MUX2X1 U429 ( .B(n580), .A(n581), .S(n1171), .Y(n579) );
  MUX2X1 U430 ( .B(n583), .A(n584), .S(n1189), .Y(n582) );
  MUX2X1 U431 ( .B(n586), .A(n587), .S(n1189), .Y(n585) );
  MUX2X1 U432 ( .B(n589), .A(n590), .S(n1189), .Y(n588) );
  MUX2X1 U433 ( .B(n592), .A(n593), .S(n1189), .Y(n591) );
  MUX2X1 U434 ( .B(n595), .A(n596), .S(n1171), .Y(n594) );
  MUX2X1 U435 ( .B(n598), .A(n599), .S(n1190), .Y(n597) );
  MUX2X1 U436 ( .B(n601), .A(n602), .S(n1190), .Y(n600) );
  MUX2X1 U437 ( .B(n604), .A(n605), .S(n1190), .Y(n603) );
  MUX2X1 U438 ( .B(n607), .A(n608), .S(n1190), .Y(n606) );
  MUX2X1 U439 ( .B(n610), .A(n611), .S(n1171), .Y(n609) );
  MUX2X1 U440 ( .B(n613), .A(n614), .S(n1190), .Y(n612) );
  MUX2X1 U441 ( .B(n616), .A(n617), .S(n1190), .Y(n615) );
  MUX2X1 U442 ( .B(n619), .A(n620), .S(n1190), .Y(n618) );
  MUX2X1 U443 ( .B(n622), .A(n623), .S(n1190), .Y(n621) );
  MUX2X1 U444 ( .B(n625), .A(n626), .S(n1171), .Y(n624) );
  MUX2X1 U445 ( .B(n628), .A(n629), .S(n1190), .Y(n627) );
  MUX2X1 U446 ( .B(n631), .A(n632), .S(n1190), .Y(n630) );
  MUX2X1 U447 ( .B(n634), .A(n635), .S(n1190), .Y(n633) );
  MUX2X1 U448 ( .B(n637), .A(n638), .S(n1190), .Y(n636) );
  MUX2X1 U449 ( .B(n640), .A(n641), .S(n1171), .Y(n639) );
  MUX2X1 U450 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n1210), .Y(n163) );
  MUX2X1 U451 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n1209), .Y(n162) );
  MUX2X1 U452 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n1209), .Y(n166) );
  MUX2X1 U453 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n1209), .Y(n165) );
  MUX2X1 U454 ( .B(n164), .A(n161), .S(n1177), .Y(n175) );
  MUX2X1 U455 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n1194), .Y(n169) );
  MUX2X1 U456 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n1194), .Y(n168) );
  MUX2X1 U457 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n1194), .Y(n172) );
  MUX2X1 U458 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n1194), .Y(n171) );
  MUX2X1 U459 ( .B(n170), .A(n167), .S(n1177), .Y(n174) );
  MUX2X1 U460 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n1194), .Y(n178) );
  MUX2X1 U461 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n1194), .Y(n177) );
  MUX2X1 U462 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n1194), .Y(n181) );
  MUX2X1 U463 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n1194), .Y(n180) );
  MUX2X1 U464 ( .B(n179), .A(n176), .S(n1177), .Y(n190) );
  MUX2X1 U465 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n1194), .Y(n184) );
  MUX2X1 U466 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n1194), .Y(n183) );
  MUX2X1 U467 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n1194), .Y(n187) );
  MUX2X1 U468 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n1194), .Y(n186) );
  MUX2X1 U469 ( .B(n185), .A(n182), .S(n1177), .Y(n189) );
  MUX2X1 U470 ( .B(n188), .A(n173), .S(n1170), .Y(n642) );
  MUX2X1 U471 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n1195), .Y(n193) );
  MUX2X1 U472 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n1195), .Y(n192) );
  MUX2X1 U473 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n1195), .Y(n196) );
  MUX2X1 U474 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n1195), .Y(n195) );
  MUX2X1 U475 ( .B(n194), .A(n191), .S(n1177), .Y(n205) );
  MUX2X1 U476 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n1195), .Y(n199) );
  MUX2X1 U477 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n1195), .Y(n198) );
  MUX2X1 U478 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n1195), .Y(n202) );
  MUX2X1 U479 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n1195), .Y(n201) );
  MUX2X1 U480 ( .B(n200), .A(n197), .S(n1177), .Y(n204) );
  MUX2X1 U481 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n1195), .Y(n208) );
  MUX2X1 U482 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n1195), .Y(n207) );
  MUX2X1 U483 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n1195), .Y(n211) );
  MUX2X1 U484 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n1195), .Y(n210) );
  MUX2X1 U485 ( .B(n209), .A(n206), .S(n1177), .Y(n221) );
  MUX2X1 U486 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n1200), .Y(n215) );
  MUX2X1 U487 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n1203), .Y(n213) );
  MUX2X1 U488 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n1200), .Y(n218) );
  MUX2X1 U489 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n1207), .Y(n217) );
  MUX2X1 U490 ( .B(n216), .A(n212), .S(n1177), .Y(n220) );
  MUX2X1 U491 ( .B(n219), .A(n203), .S(n1170), .Y(n643) );
  MUX2X1 U492 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n1206), .Y(n224) );
  MUX2X1 U493 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n1199), .Y(n223) );
  MUX2X1 U494 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n1205), .Y(n227) );
  MUX2X1 U495 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n1202), .Y(n226) );
  MUX2X1 U496 ( .B(n225), .A(n222), .S(n1177), .Y(n236) );
  MUX2X1 U497 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n1207), .Y(n230) );
  MUX2X1 U498 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n1208), .Y(n229) );
  MUX2X1 U499 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n1204), .Y(n233) );
  MUX2X1 U500 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n1209), .Y(n232) );
  MUX2X1 U501 ( .B(n231), .A(n228), .S(n1177), .Y(n235) );
  MUX2X1 U502 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n1196), .Y(n239) );
  MUX2X1 U503 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n1196), .Y(n238) );
  MUX2X1 U504 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n1196), .Y(n242) );
  MUX2X1 U505 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n1196), .Y(n241) );
  MUX2X1 U506 ( .B(n240), .A(n237), .S(n1177), .Y(n251) );
  MUX2X1 U507 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n1196), .Y(n245) );
  MUX2X1 U508 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n1196), .Y(n244) );
  MUX2X1 U509 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n1196), .Y(n248) );
  MUX2X1 U510 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n1196), .Y(n247) );
  MUX2X1 U511 ( .B(n246), .A(n243), .S(n1177), .Y(n250) );
  MUX2X1 U512 ( .B(n249), .A(n234), .S(n1170), .Y(n644) );
  MUX2X1 U513 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n1196), .Y(n254) );
  MUX2X1 U514 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n1196), .Y(n253) );
  MUX2X1 U515 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n1196), .Y(n257) );
  MUX2X1 U516 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n1196), .Y(n256) );
  MUX2X1 U517 ( .B(n255), .A(n252), .S(n1176), .Y(n266) );
  MUX2X1 U518 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n1197), .Y(n260) );
  MUX2X1 U519 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n1197), .Y(n259) );
  MUX2X1 U520 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n1197), .Y(n263) );
  MUX2X1 U521 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n1197), .Y(n262) );
  MUX2X1 U522 ( .B(n261), .A(n258), .S(n1176), .Y(n265) );
  MUX2X1 U523 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n1197), .Y(n269) );
  MUX2X1 U524 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n1197), .Y(n268) );
  MUX2X1 U525 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n1197), .Y(n272) );
  MUX2X1 U526 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n1197), .Y(n271) );
  MUX2X1 U527 ( .B(n270), .A(n267), .S(n1176), .Y(n281) );
  MUX2X1 U528 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n1197), .Y(n275) );
  MUX2X1 U529 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n1197), .Y(n274) );
  MUX2X1 U530 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n1197), .Y(n278) );
  MUX2X1 U531 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n1197), .Y(n277) );
  MUX2X1 U532 ( .B(n276), .A(n273), .S(n1176), .Y(n280) );
  MUX2X1 U533 ( .B(n279), .A(n264), .S(n1170), .Y(n645) );
  MUX2X1 U534 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n1198), .Y(n284) );
  MUX2X1 U535 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n1198), .Y(n283) );
  MUX2X1 U536 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n1198), .Y(n287) );
  MUX2X1 U537 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n1198), .Y(n286) );
  MUX2X1 U538 ( .B(n285), .A(n282), .S(n1176), .Y(n296) );
  MUX2X1 U539 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n1198), .Y(n290) );
  MUX2X1 U540 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n1198), .Y(n289) );
  MUX2X1 U541 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n1198), .Y(n293) );
  MUX2X1 U542 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n1198), .Y(n292) );
  MUX2X1 U543 ( .B(n291), .A(n288), .S(n1176), .Y(n295) );
  MUX2X1 U544 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n1198), .Y(n299) );
  MUX2X1 U545 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n1198), .Y(n298) );
  MUX2X1 U546 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n1198), .Y(n302) );
  MUX2X1 U547 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n1198), .Y(n301) );
  MUX2X1 U548 ( .B(n300), .A(n297), .S(n1176), .Y(n311) );
  MUX2X1 U549 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n1199), .Y(n305) );
  MUX2X1 U550 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n1199), .Y(n304) );
  MUX2X1 U551 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n1199), .Y(n308) );
  MUX2X1 U552 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n1199), .Y(n307) );
  MUX2X1 U553 ( .B(n306), .A(n303), .S(n1176), .Y(n310) );
  MUX2X1 U554 ( .B(n309), .A(n294), .S(n1170), .Y(n646) );
  MUX2X1 U555 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n1199), .Y(n314) );
  MUX2X1 U556 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n1199), .Y(n313) );
  MUX2X1 U557 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n1199), .Y(n317) );
  MUX2X1 U558 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n1199), .Y(n316) );
  MUX2X1 U559 ( .B(n315), .A(n312), .S(n1176), .Y(n326) );
  MUX2X1 U560 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n1199), .Y(n320) );
  MUX2X1 U561 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n1199), .Y(n319) );
  MUX2X1 U562 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n1199), .Y(n323) );
  MUX2X1 U563 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n1199), .Y(n322) );
  MUX2X1 U564 ( .B(n321), .A(n318), .S(n1176), .Y(n325) );
  MUX2X1 U565 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n1200), .Y(n329) );
  MUX2X1 U566 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n1200), .Y(n328) );
  MUX2X1 U567 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n1200), .Y(n332) );
  MUX2X1 U568 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n1200), .Y(n331) );
  MUX2X1 U569 ( .B(n330), .A(n327), .S(n1176), .Y(n341) );
  MUX2X1 U570 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n1200), .Y(n335) );
  MUX2X1 U571 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n1200), .Y(n334) );
  MUX2X1 U572 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n1200), .Y(n338) );
  MUX2X1 U573 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n1200), .Y(n337) );
  MUX2X1 U574 ( .B(n336), .A(n333), .S(n1176), .Y(n340) );
  MUX2X1 U575 ( .B(n339), .A(n324), .S(n1170), .Y(n647) );
  MUX2X1 U576 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n1200), .Y(n344) );
  MUX2X1 U577 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n1200), .Y(n343) );
  MUX2X1 U578 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n1200), .Y(n347) );
  MUX2X1 U579 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n1200), .Y(n346) );
  MUX2X1 U580 ( .B(n345), .A(n342), .S(n1177), .Y(n356) );
  MUX2X1 U581 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n1199), .Y(n350) );
  MUX2X1 U582 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n1207), .Y(n349) );
  MUX2X1 U583 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n1208), .Y(n353) );
  MUX2X1 U584 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n1208), .Y(n352) );
  MUX2X1 U585 ( .B(n351), .A(n348), .S(n1176), .Y(n355) );
  MUX2X1 U586 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n1207), .Y(n359) );
  MUX2X1 U587 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n1208), .Y(n358) );
  MUX2X1 U588 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n1201), .Y(n362) );
  MUX2X1 U589 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n1202), .Y(n361) );
  MUX2X1 U590 ( .B(n360), .A(n357), .S(n1176), .Y(n371) );
  MUX2X1 U591 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n1199), .Y(n365) );
  MUX2X1 U592 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n1199), .Y(n364) );
  MUX2X1 U593 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n1204), .Y(n368) );
  MUX2X1 U594 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n1198), .Y(n367) );
  MUX2X1 U595 ( .B(n366), .A(n363), .S(n1176), .Y(n370) );
  MUX2X1 U596 ( .B(n369), .A(n354), .S(n1170), .Y(n648) );
  MUX2X1 U597 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n1208), .Y(n374) );
  MUX2X1 U598 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n1200), .Y(n373) );
  MUX2X1 U599 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n1208), .Y(n377) );
  MUX2X1 U600 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n1200), .Y(n376) );
  MUX2X1 U601 ( .B(n375), .A(n372), .S(n1177), .Y(n386) );
  MUX2X1 U602 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n1199), .Y(n380) );
  MUX2X1 U603 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n1207), .Y(n379) );
  MUX2X1 U604 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n1208), .Y(n383) );
  MUX2X1 U605 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n1207), .Y(n382) );
  MUX2X1 U606 ( .B(n381), .A(n378), .S(n1176), .Y(n385) );
  MUX2X1 U607 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n1199), .Y(n389) );
  MUX2X1 U608 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n1199), .Y(n388) );
  MUX2X1 U609 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n1198), .Y(n392) );
  MUX2X1 U610 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n1200), .Y(n391) );
  MUX2X1 U611 ( .B(n390), .A(n387), .S(n1177), .Y(n401) );
  MUX2X1 U612 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n1200), .Y(n395) );
  MUX2X1 U613 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n1200), .Y(n394) );
  MUX2X1 U614 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n1198), .Y(n398) );
  MUX2X1 U615 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n1200), .Y(n397) );
  MUX2X1 U616 ( .B(n396), .A(n393), .S(n1176), .Y(n400) );
  MUX2X1 U617 ( .B(n399), .A(n384), .S(n1170), .Y(n649) );
  MUX2X1 U618 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n1200), .Y(n404) );
  MUX2X1 U619 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n1198), .Y(n403) );
  MUX2X1 U620 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n1198), .Y(n407) );
  MUX2X1 U621 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n1198), .Y(n406) );
  MUX2X1 U622 ( .B(n405), .A(n402), .S(n1176), .Y(n416) );
  MUX2X1 U623 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n1200), .Y(n410) );
  MUX2X1 U624 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n1198), .Y(n409) );
  MUX2X1 U625 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n1198), .Y(n413) );
  MUX2X1 U626 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n1198), .Y(n412) );
  MUX2X1 U627 ( .B(n411), .A(n408), .S(n1177), .Y(n415) );
  MUX2X1 U628 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n1201), .Y(n419) );
  MUX2X1 U629 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n1201), .Y(n418) );
  MUX2X1 U630 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n1201), .Y(n422) );
  MUX2X1 U631 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n1201), .Y(n421) );
  MUX2X1 U632 ( .B(n420), .A(n417), .S(n1176), .Y(n431) );
  MUX2X1 U633 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n1201), .Y(n425) );
  MUX2X1 U634 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n1201), .Y(n424) );
  MUX2X1 U635 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n1201), .Y(n428) );
  MUX2X1 U636 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n1201), .Y(n427) );
  MUX2X1 U637 ( .B(n426), .A(n423), .S(n1177), .Y(n430) );
  MUX2X1 U638 ( .B(n429), .A(n414), .S(n1170), .Y(n650) );
  MUX2X1 U639 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n1201), .Y(n434) );
  MUX2X1 U640 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n1201), .Y(n433) );
  MUX2X1 U641 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n1201), .Y(n437) );
  MUX2X1 U642 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n1201), .Y(n436) );
  MUX2X1 U643 ( .B(n435), .A(n432), .S(n1175), .Y(n446) );
  MUX2X1 U644 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n1202), .Y(n440) );
  MUX2X1 U645 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n1202), .Y(n439) );
  MUX2X1 U646 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n1202), .Y(n443) );
  MUX2X1 U647 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n1202), .Y(n442) );
  MUX2X1 U648 ( .B(n441), .A(n438), .S(n1175), .Y(n445) );
  MUX2X1 U649 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n1202), .Y(n449) );
  MUX2X1 U650 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n1202), .Y(n448) );
  MUX2X1 U651 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n1202), .Y(n452) );
  MUX2X1 U652 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n1202), .Y(n451) );
  MUX2X1 U653 ( .B(n450), .A(n447), .S(n1175), .Y(n461) );
  MUX2X1 U654 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n1202), .Y(n455) );
  MUX2X1 U655 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n1202), .Y(n454) );
  MUX2X1 U656 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n1202), .Y(n458) );
  MUX2X1 U657 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n1202), .Y(n457) );
  MUX2X1 U658 ( .B(n456), .A(n453), .S(n1175), .Y(n460) );
  MUX2X1 U659 ( .B(n459), .A(n444), .S(n1170), .Y(n1163) );
  MUX2X1 U660 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n1203), .Y(n464) );
  MUX2X1 U661 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n1203), .Y(n463) );
  MUX2X1 U662 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n1203), .Y(n467) );
  MUX2X1 U663 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n1203), .Y(n466) );
  MUX2X1 U664 ( .B(n465), .A(n462), .S(n1175), .Y(n476) );
  MUX2X1 U665 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n1203), .Y(n470) );
  MUX2X1 U666 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n1203), .Y(n469) );
  MUX2X1 U667 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n1203), .Y(n473) );
  MUX2X1 U668 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n1203), .Y(n472) );
  MUX2X1 U669 ( .B(n471), .A(n468), .S(n1175), .Y(n475) );
  MUX2X1 U670 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n1203), .Y(n479) );
  MUX2X1 U671 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n1203), .Y(n478) );
  MUX2X1 U672 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n1203), .Y(n482) );
  MUX2X1 U673 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n1203), .Y(n481) );
  MUX2X1 U674 ( .B(n480), .A(n477), .S(n1175), .Y(n491) );
  MUX2X1 U675 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n1204), .Y(n485) );
  MUX2X1 U676 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n1204), .Y(n484) );
  MUX2X1 U677 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n1204), .Y(n488) );
  MUX2X1 U678 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n1204), .Y(n487) );
  MUX2X1 U679 ( .B(n486), .A(n483), .S(n1175), .Y(n490) );
  MUX2X1 U680 ( .B(n489), .A(n474), .S(n1170), .Y(n1164) );
  MUX2X1 U681 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n1204), .Y(n494) );
  MUX2X1 U682 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n1204), .Y(n493) );
  MUX2X1 U683 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n1204), .Y(n497) );
  MUX2X1 U684 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n1204), .Y(n496) );
  MUX2X1 U685 ( .B(n495), .A(n492), .S(n1175), .Y(n506) );
  MUX2X1 U686 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n1204), .Y(n500) );
  MUX2X1 U687 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n1204), .Y(n499) );
  MUX2X1 U688 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n1204), .Y(n503) );
  MUX2X1 U689 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n1204), .Y(n502) );
  MUX2X1 U690 ( .B(n501), .A(n498), .S(n1175), .Y(n505) );
  MUX2X1 U691 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n1205), .Y(n509) );
  MUX2X1 U692 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n1205), .Y(n508) );
  MUX2X1 U693 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n1205), .Y(n512) );
  MUX2X1 U694 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n1205), .Y(n511) );
  MUX2X1 U695 ( .B(n510), .A(n507), .S(n1175), .Y(n521) );
  MUX2X1 U696 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n1205), .Y(n515) );
  MUX2X1 U697 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n1205), .Y(n514) );
  MUX2X1 U698 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n1205), .Y(n518) );
  MUX2X1 U699 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n1205), .Y(n517) );
  MUX2X1 U700 ( .B(n516), .A(n513), .S(n1175), .Y(n520) );
  MUX2X1 U701 ( .B(n519), .A(n504), .S(n1170), .Y(n1165) );
  MUX2X1 U702 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n1205), .Y(n524) );
  MUX2X1 U703 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n1205), .Y(n523) );
  MUX2X1 U704 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n1205), .Y(n527) );
  MUX2X1 U705 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n1205), .Y(n526) );
  MUX2X1 U706 ( .B(n525), .A(n522), .S(n1174), .Y(n536) );
  MUX2X1 U707 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n1206), .Y(n530) );
  MUX2X1 U708 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n1206), .Y(n529) );
  MUX2X1 U709 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n1206), .Y(n533) );
  MUX2X1 U710 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n1206), .Y(n532) );
  MUX2X1 U711 ( .B(n531), .A(n528), .S(n1174), .Y(n535) );
  MUX2X1 U712 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n1206), .Y(n539) );
  MUX2X1 U713 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n1206), .Y(n538) );
  MUX2X1 U714 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n1206), .Y(n542) );
  MUX2X1 U715 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n1206), .Y(n541) );
  MUX2X1 U716 ( .B(n540), .A(n537), .S(n1174), .Y(n551) );
  MUX2X1 U717 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n1206), .Y(n545) );
  MUX2X1 U718 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n1206), .Y(n544) );
  MUX2X1 U719 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n1206), .Y(n548) );
  MUX2X1 U720 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n1206), .Y(n547) );
  MUX2X1 U721 ( .B(n546), .A(n543), .S(n1174), .Y(n550) );
  MUX2X1 U722 ( .B(n549), .A(n534), .S(n1170), .Y(n1166) );
  MUX2X1 U723 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n1207), .Y(n554) );
  MUX2X1 U724 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n1207), .Y(n553) );
  MUX2X1 U725 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n1207), .Y(n557) );
  MUX2X1 U726 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n1207), .Y(n556) );
  MUX2X1 U727 ( .B(n555), .A(n552), .S(n1174), .Y(n566) );
  MUX2X1 U728 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n1207), .Y(n560) );
  MUX2X1 U729 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n1207), .Y(n559) );
  MUX2X1 U730 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n1207), .Y(n563) );
  MUX2X1 U731 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n1207), .Y(n562) );
  MUX2X1 U732 ( .B(n561), .A(n558), .S(n1174), .Y(n565) );
  MUX2X1 U733 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n1207), .Y(n569) );
  MUX2X1 U734 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n1207), .Y(n568) );
  MUX2X1 U735 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n1207), .Y(n572) );
  MUX2X1 U736 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n1207), .Y(n571) );
  MUX2X1 U737 ( .B(n570), .A(n567), .S(n1174), .Y(n581) );
  MUX2X1 U738 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n1208), .Y(n575) );
  MUX2X1 U739 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n1208), .Y(n574) );
  MUX2X1 U740 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n1208), .Y(n578) );
  MUX2X1 U741 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n1208), .Y(n577) );
  MUX2X1 U742 ( .B(n576), .A(n573), .S(n1174), .Y(n580) );
  MUX2X1 U743 ( .B(n579), .A(n564), .S(n1170), .Y(n1167) );
  MUX2X1 U744 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n1208), .Y(n584) );
  MUX2X1 U745 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n1208), .Y(n583) );
  MUX2X1 U746 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n1208), .Y(n587) );
  MUX2X1 U747 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n1208), .Y(n586) );
  MUX2X1 U748 ( .B(n585), .A(n582), .S(n1174), .Y(n596) );
  MUX2X1 U749 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n1208), .Y(n590) );
  MUX2X1 U750 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n1208), .Y(n589) );
  MUX2X1 U751 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n1208), .Y(n593) );
  MUX2X1 U752 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n1208), .Y(n592) );
  MUX2X1 U753 ( .B(n591), .A(n588), .S(n1174), .Y(n595) );
  MUX2X1 U754 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n1209), .Y(n599) );
  MUX2X1 U755 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n1209), .Y(n598) );
  MUX2X1 U756 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n1209), .Y(n602) );
  MUX2X1 U757 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n1209), .Y(n601) );
  MUX2X1 U758 ( .B(n600), .A(n597), .S(n1174), .Y(n611) );
  MUX2X1 U759 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n1209), .Y(n605) );
  MUX2X1 U760 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n1209), .Y(n604) );
  MUX2X1 U761 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n1209), .Y(n608) );
  MUX2X1 U762 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n1209), .Y(n607) );
  MUX2X1 U763 ( .B(n606), .A(n603), .S(n1174), .Y(n610) );
  MUX2X1 U764 ( .B(n609), .A(n594), .S(n1170), .Y(n1168) );
  MUX2X1 U765 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n1209), .Y(n614) );
  MUX2X1 U766 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n1209), .Y(n613) );
  MUX2X1 U767 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n1209), .Y(n617) );
  MUX2X1 U768 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n1209), .Y(n616) );
  MUX2X1 U769 ( .B(n615), .A(n612), .S(n1175), .Y(n626) );
  MUX2X1 U770 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n1210), .Y(n620) );
  MUX2X1 U771 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n1210), .Y(n619) );
  MUX2X1 U772 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n1210), .Y(n623) );
  MUX2X1 U773 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n1210), .Y(n622) );
  MUX2X1 U774 ( .B(n621), .A(n618), .S(n1174), .Y(n625) );
  MUX2X1 U775 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n1210), .Y(n629) );
  MUX2X1 U776 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n1210), .Y(n628) );
  MUX2X1 U777 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n1210), .Y(n632) );
  MUX2X1 U778 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n1210), .Y(n631) );
  MUX2X1 U779 ( .B(n630), .A(n627), .S(n1175), .Y(n641) );
  MUX2X1 U780 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n1210), .Y(n635) );
  MUX2X1 U781 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n1210), .Y(n634) );
  MUX2X1 U782 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n1210), .Y(n638) );
  MUX2X1 U783 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n1210), .Y(n637) );
  MUX2X1 U784 ( .B(n636), .A(n633), .S(n1174), .Y(n640) );
  MUX2X1 U785 ( .B(n639), .A(n624), .S(n1170), .Y(n1169) );
  INVX1 U786 ( .A(N12), .Y(n1299) );
  INVX1 U787 ( .A(N11), .Y(n1297) );
  INVX8 U788 ( .A(n1269), .Y(n1266) );
  INVX8 U789 ( .A(n1269), .Y(n1267) );
  INVX8 U790 ( .A(n1269), .Y(n1268) );
  INVX8 U791 ( .A(n59), .Y(n1269) );
  INVX8 U792 ( .A(n73), .Y(n1270) );
  INVX8 U793 ( .A(n74), .Y(n1271) );
  INVX8 U794 ( .A(n74), .Y(n1272) );
  INVX8 U795 ( .A(n75), .Y(n1273) );
  INVX8 U796 ( .A(n76), .Y(n1274) );
  INVX8 U797 ( .A(n77), .Y(n1275) );
  INVX8 U798 ( .A(n78), .Y(n1276) );
  INVX8 U799 ( .A(n78), .Y(n1277) );
  INVX8 U800 ( .A(n79), .Y(n1278) );
  INVX8 U801 ( .A(n80), .Y(n1279) );
  INVX8 U802 ( .A(n81), .Y(n1280) );
  INVX8 U803 ( .A(n82), .Y(n1281) );
  INVX8 U804 ( .A(n82), .Y(n1282) );
  INVX8 U805 ( .A(n83), .Y(n1283) );
  INVX8 U806 ( .A(n84), .Y(n1284) );
  INVX8 U807 ( .A(n84), .Y(n1285) );
  INVX8 U808 ( .A(n85), .Y(n1286) );
  INVX8 U809 ( .A(n85), .Y(n1287) );
  INVX8 U810 ( .A(n86), .Y(n1288) );
  INVX8 U811 ( .A(n86), .Y(n1289) );
  INVX8 U812 ( .A(n87), .Y(n1290) );
  INVX8 U813 ( .A(n87), .Y(n1291) );
  INVX8 U814 ( .A(n88), .Y(n1292) );
  INVX8 U815 ( .A(n88), .Y(n1293) );
  OR2X2 U816 ( .A(write), .B(rst), .Y(n1304) );
  AND2X2 U817 ( .A(N32), .B(n1305), .Y(\data_out<0> ) );
  AND2X2 U818 ( .A(n1), .B(N31), .Y(\data_out<1> ) );
  AND2X2 U819 ( .A(N30), .B(n1305), .Y(\data_out<2> ) );
  AND2X2 U820 ( .A(n1), .B(N29), .Y(\data_out<3> ) );
  AND2X2 U821 ( .A(N28), .B(n1305), .Y(\data_out<4> ) );
  AND2X2 U822 ( .A(N27), .B(n1305), .Y(\data_out<5> ) );
  AND2X2 U823 ( .A(N26), .B(n1), .Y(\data_out<6> ) );
  AND2X2 U824 ( .A(N25), .B(n1305), .Y(\data_out<7> ) );
  AND2X2 U825 ( .A(N24), .B(n1), .Y(\data_out<8> ) );
  AND2X2 U826 ( .A(N23), .B(n1), .Y(\data_out<9> ) );
  AND2X2 U827 ( .A(N22), .B(n1305), .Y(\data_out<10> ) );
  AND2X2 U828 ( .A(n1), .B(N21), .Y(\data_out<11> ) );
  AND2X2 U829 ( .A(N20), .B(n1305), .Y(\data_out<12> ) );
  AND2X2 U830 ( .A(N19), .B(n1), .Y(\data_out<13> ) );
  AND2X2 U831 ( .A(N18), .B(n1), .Y(\data_out<14> ) );
  AND2X2 U832 ( .A(N17), .B(n1305), .Y(\data_out<15> ) );
  NAND2X1 U833 ( .A(\mem<31><0> ), .B(n1212), .Y(n1306) );
  OAI21X1 U834 ( .A(n94), .B(n1270), .C(n1306), .Y(n2344) );
  NAND2X1 U835 ( .A(\mem<31><1> ), .B(n1212), .Y(n1307) );
  OAI21X1 U836 ( .A(n1272), .B(n94), .C(n1307), .Y(n2343) );
  NAND2X1 U837 ( .A(\mem<31><2> ), .B(n1212), .Y(n1308) );
  OAI21X1 U838 ( .A(n1273), .B(n94), .C(n1308), .Y(n2342) );
  NAND2X1 U839 ( .A(\mem<31><3> ), .B(n1212), .Y(n1309) );
  OAI21X1 U840 ( .A(n1274), .B(n94), .C(n1309), .Y(n2341) );
  NAND2X1 U841 ( .A(\mem<31><4> ), .B(n1212), .Y(n1310) );
  OAI21X1 U842 ( .A(n1275), .B(n94), .C(n1310), .Y(n2340) );
  NAND2X1 U843 ( .A(\mem<31><5> ), .B(n1212), .Y(n1311) );
  OAI21X1 U844 ( .A(n1277), .B(n94), .C(n1311), .Y(n2339) );
  NAND2X1 U845 ( .A(\mem<31><6> ), .B(n1212), .Y(n1312) );
  OAI21X1 U846 ( .A(n1278), .B(n94), .C(n1312), .Y(n2338) );
  NAND2X1 U847 ( .A(\mem<31><7> ), .B(n1212), .Y(n1313) );
  OAI21X1 U848 ( .A(n1279), .B(n94), .C(n1313), .Y(n2337) );
  NAND2X1 U849 ( .A(\mem<31><8> ), .B(n1213), .Y(n1314) );
  OAI21X1 U850 ( .A(n1280), .B(n94), .C(n1314), .Y(n2336) );
  NAND2X1 U851 ( .A(\mem<31><9> ), .B(n1213), .Y(n1315) );
  OAI21X1 U852 ( .A(n1282), .B(n94), .C(n1315), .Y(n2335) );
  NAND2X1 U853 ( .A(\mem<31><10> ), .B(n1213), .Y(n1316) );
  OAI21X1 U854 ( .A(n1283), .B(n94), .C(n1316), .Y(n2334) );
  NAND2X1 U855 ( .A(\mem<31><11> ), .B(n1213), .Y(n1317) );
  OAI21X1 U856 ( .A(n1285), .B(n94), .C(n1317), .Y(n2333) );
  NAND2X1 U857 ( .A(\mem<31><12> ), .B(n1213), .Y(n1318) );
  OAI21X1 U858 ( .A(n1287), .B(n94), .C(n1318), .Y(n2332) );
  NAND2X1 U859 ( .A(\mem<31><13> ), .B(n1213), .Y(n1319) );
  OAI21X1 U860 ( .A(n1289), .B(n94), .C(n1319), .Y(n2331) );
  NAND2X1 U861 ( .A(\mem<31><14> ), .B(n1213), .Y(n1320) );
  OAI21X1 U862 ( .A(n1291), .B(n94), .C(n1320), .Y(n2330) );
  NAND2X1 U863 ( .A(\mem<31><15> ), .B(n1213), .Y(n1321) );
  OAI21X1 U864 ( .A(n1293), .B(n94), .C(n1321), .Y(n2329) );
  NAND2X1 U865 ( .A(\mem<30><0> ), .B(n1214), .Y(n1322) );
  OAI21X1 U866 ( .A(n96), .B(n1270), .C(n1322), .Y(n2328) );
  NAND2X1 U867 ( .A(\mem<30><1> ), .B(n1214), .Y(n1323) );
  OAI21X1 U868 ( .A(n96), .B(n1272), .C(n1323), .Y(n2327) );
  NAND2X1 U869 ( .A(\mem<30><2> ), .B(n1214), .Y(n1324) );
  OAI21X1 U870 ( .A(n96), .B(n1273), .C(n1324), .Y(n2326) );
  NAND2X1 U871 ( .A(\mem<30><3> ), .B(n1214), .Y(n1325) );
  OAI21X1 U872 ( .A(n96), .B(n1274), .C(n1325), .Y(n2325) );
  NAND2X1 U873 ( .A(\mem<30><4> ), .B(n1214), .Y(n1326) );
  OAI21X1 U874 ( .A(n96), .B(n1275), .C(n1326), .Y(n2324) );
  NAND2X1 U875 ( .A(\mem<30><5> ), .B(n1214), .Y(n1327) );
  OAI21X1 U876 ( .A(n96), .B(n1277), .C(n1327), .Y(n2323) );
  NAND2X1 U877 ( .A(\mem<30><6> ), .B(n1214), .Y(n1328) );
  OAI21X1 U878 ( .A(n96), .B(n1278), .C(n1328), .Y(n2322) );
  NAND2X1 U879 ( .A(\mem<30><7> ), .B(n1214), .Y(n1329) );
  OAI21X1 U880 ( .A(n96), .B(n1279), .C(n1329), .Y(n2321) );
  NAND2X1 U881 ( .A(\mem<30><8> ), .B(n1215), .Y(n1330) );
  OAI21X1 U882 ( .A(n96), .B(n1280), .C(n1330), .Y(n2320) );
  NAND2X1 U883 ( .A(\mem<30><9> ), .B(n1215), .Y(n1331) );
  OAI21X1 U884 ( .A(n96), .B(n1281), .C(n1331), .Y(n2319) );
  NAND2X1 U885 ( .A(\mem<30><10> ), .B(n1215), .Y(n1332) );
  OAI21X1 U886 ( .A(n96), .B(n1283), .C(n1332), .Y(n2318) );
  NAND2X1 U887 ( .A(\mem<30><11> ), .B(n1215), .Y(n1333) );
  OAI21X1 U888 ( .A(n96), .B(n1284), .C(n1333), .Y(n2317) );
  NAND2X1 U889 ( .A(\mem<30><12> ), .B(n1215), .Y(n1334) );
  OAI21X1 U890 ( .A(n96), .B(n1286), .C(n1334), .Y(n2316) );
  NAND2X1 U891 ( .A(\mem<30><13> ), .B(n1215), .Y(n1335) );
  OAI21X1 U892 ( .A(n96), .B(n1288), .C(n1335), .Y(n2315) );
  NAND2X1 U893 ( .A(\mem<30><14> ), .B(n1215), .Y(n1336) );
  OAI21X1 U894 ( .A(n96), .B(n1290), .C(n1336), .Y(n2314) );
  NAND2X1 U895 ( .A(\mem<30><15> ), .B(n1215), .Y(n1337) );
  OAI21X1 U896 ( .A(n96), .B(n1292), .C(n1337), .Y(n2313) );
  NAND3X1 U897 ( .A(N10), .B(n1298), .C(n1297), .Y(n1338) );
  NAND2X1 U898 ( .A(\mem<29><0> ), .B(n1216), .Y(n1339) );
  OAI21X1 U899 ( .A(n98), .B(n1270), .C(n1339), .Y(n2312) );
  NAND2X1 U900 ( .A(\mem<29><1> ), .B(n1216), .Y(n1340) );
  OAI21X1 U901 ( .A(n98), .B(n1271), .C(n1340), .Y(n2311) );
  NAND2X1 U902 ( .A(\mem<29><2> ), .B(n1216), .Y(n1341) );
  OAI21X1 U903 ( .A(n98), .B(n1273), .C(n1341), .Y(n2310) );
  NAND2X1 U904 ( .A(\mem<29><3> ), .B(n1216), .Y(n1342) );
  OAI21X1 U905 ( .A(n98), .B(n1274), .C(n1342), .Y(n2309) );
  NAND2X1 U906 ( .A(\mem<29><4> ), .B(n1216), .Y(n1343) );
  OAI21X1 U907 ( .A(n98), .B(n1275), .C(n1343), .Y(n2308) );
  NAND2X1 U908 ( .A(\mem<29><5> ), .B(n1216), .Y(n1344) );
  OAI21X1 U909 ( .A(n98), .B(n1276), .C(n1344), .Y(n2307) );
  NAND2X1 U910 ( .A(\mem<29><6> ), .B(n1216), .Y(n1345) );
  OAI21X1 U911 ( .A(n98), .B(n1278), .C(n1345), .Y(n2306) );
  NAND2X1 U912 ( .A(\mem<29><7> ), .B(n1216), .Y(n1346) );
  OAI21X1 U913 ( .A(n98), .B(n1279), .C(n1346), .Y(n2305) );
  NAND2X1 U914 ( .A(\mem<29><8> ), .B(n1217), .Y(n1347) );
  OAI21X1 U915 ( .A(n98), .B(n1280), .C(n1347), .Y(n2304) );
  NAND2X1 U916 ( .A(\mem<29><9> ), .B(n1217), .Y(n1348) );
  OAI21X1 U917 ( .A(n98), .B(n1282), .C(n1348), .Y(n2303) );
  NAND2X1 U918 ( .A(\mem<29><10> ), .B(n1217), .Y(n1349) );
  OAI21X1 U919 ( .A(n98), .B(n1283), .C(n1349), .Y(n2302) );
  NAND2X1 U920 ( .A(\mem<29><11> ), .B(n1217), .Y(n1350) );
  OAI21X1 U921 ( .A(n98), .B(n1285), .C(n1350), .Y(n2301) );
  NAND2X1 U922 ( .A(\mem<29><12> ), .B(n1217), .Y(n1351) );
  OAI21X1 U923 ( .A(n98), .B(n1287), .C(n1351), .Y(n2300) );
  NAND2X1 U924 ( .A(\mem<29><13> ), .B(n1217), .Y(n1352) );
  OAI21X1 U925 ( .A(n98), .B(n1289), .C(n1352), .Y(n2299) );
  NAND2X1 U926 ( .A(\mem<29><14> ), .B(n1217), .Y(n1353) );
  OAI21X1 U927 ( .A(n98), .B(n1291), .C(n1353), .Y(n2298) );
  NAND2X1 U928 ( .A(\mem<29><15> ), .B(n1217), .Y(n1354) );
  OAI21X1 U929 ( .A(n98), .B(n1293), .C(n1354), .Y(n2297) );
  NAND3X1 U930 ( .A(n1298), .B(n1297), .C(n1295), .Y(n1355) );
  NAND2X1 U931 ( .A(\mem<28><0> ), .B(n1218), .Y(n1356) );
  OAI21X1 U932 ( .A(n100), .B(n1270), .C(n1356), .Y(n2296) );
  NAND2X1 U933 ( .A(\mem<28><1> ), .B(n1218), .Y(n1357) );
  OAI21X1 U934 ( .A(n100), .B(n1272), .C(n1357), .Y(n2295) );
  NAND2X1 U935 ( .A(\mem<28><2> ), .B(n1218), .Y(n1358) );
  OAI21X1 U936 ( .A(n100), .B(n1273), .C(n1358), .Y(n2294) );
  NAND2X1 U937 ( .A(\mem<28><3> ), .B(n1218), .Y(n1359) );
  OAI21X1 U938 ( .A(n100), .B(n1274), .C(n1359), .Y(n2293) );
  NAND2X1 U939 ( .A(\mem<28><4> ), .B(n1218), .Y(n1360) );
  OAI21X1 U940 ( .A(n100), .B(n1275), .C(n1360), .Y(n2292) );
  NAND2X1 U941 ( .A(\mem<28><5> ), .B(n1218), .Y(n1361) );
  OAI21X1 U942 ( .A(n100), .B(n1277), .C(n1361), .Y(n2291) );
  NAND2X1 U943 ( .A(\mem<28><6> ), .B(n1218), .Y(n1362) );
  OAI21X1 U944 ( .A(n100), .B(n1278), .C(n1362), .Y(n2290) );
  NAND2X1 U945 ( .A(\mem<28><7> ), .B(n1218), .Y(n1363) );
  OAI21X1 U946 ( .A(n100), .B(n1279), .C(n1363), .Y(n2289) );
  NAND2X1 U947 ( .A(\mem<28><8> ), .B(n1219), .Y(n1364) );
  OAI21X1 U948 ( .A(n100), .B(n1280), .C(n1364), .Y(n2288) );
  NAND2X1 U949 ( .A(\mem<28><9> ), .B(n1219), .Y(n1365) );
  OAI21X1 U950 ( .A(n100), .B(n1281), .C(n1365), .Y(n2287) );
  NAND2X1 U951 ( .A(\mem<28><10> ), .B(n1219), .Y(n1366) );
  OAI21X1 U952 ( .A(n100), .B(n1283), .C(n1366), .Y(n2286) );
  NAND2X1 U953 ( .A(\mem<28><11> ), .B(n1219), .Y(n1367) );
  OAI21X1 U954 ( .A(n100), .B(n1284), .C(n1367), .Y(n2285) );
  NAND2X1 U955 ( .A(\mem<28><12> ), .B(n1219), .Y(n1368) );
  OAI21X1 U956 ( .A(n100), .B(n1286), .C(n1368), .Y(n2284) );
  NAND2X1 U957 ( .A(\mem<28><13> ), .B(n1219), .Y(n1369) );
  OAI21X1 U958 ( .A(n100), .B(n1288), .C(n1369), .Y(n2283) );
  NAND2X1 U959 ( .A(\mem<28><14> ), .B(n1219), .Y(n1370) );
  OAI21X1 U960 ( .A(n100), .B(n1290), .C(n1370), .Y(n2282) );
  NAND2X1 U961 ( .A(\mem<28><15> ), .B(n1219), .Y(n1371) );
  OAI21X1 U962 ( .A(n100), .B(n1292), .C(n1371), .Y(n2281) );
  NAND3X1 U963 ( .A(N10), .B(n1296), .C(n1299), .Y(n1372) );
  NAND2X1 U964 ( .A(\mem<27><0> ), .B(n1220), .Y(n1373) );
  OAI21X1 U965 ( .A(n102), .B(n1270), .C(n1373), .Y(n2280) );
  NAND2X1 U966 ( .A(\mem<27><1> ), .B(n1220), .Y(n1374) );
  OAI21X1 U967 ( .A(n102), .B(n1271), .C(n1374), .Y(n2279) );
  NAND2X1 U968 ( .A(\mem<27><2> ), .B(n1220), .Y(n1375) );
  OAI21X1 U969 ( .A(n102), .B(n1273), .C(n1375), .Y(n2278) );
  NAND2X1 U970 ( .A(\mem<27><3> ), .B(n1220), .Y(n1376) );
  OAI21X1 U971 ( .A(n102), .B(n1274), .C(n1376), .Y(n2277) );
  NAND2X1 U972 ( .A(\mem<27><4> ), .B(n1220), .Y(n1377) );
  OAI21X1 U973 ( .A(n102), .B(n1275), .C(n1377), .Y(n2276) );
  NAND2X1 U974 ( .A(\mem<27><5> ), .B(n1220), .Y(n1378) );
  OAI21X1 U975 ( .A(n102), .B(n1276), .C(n1378), .Y(n2275) );
  NAND2X1 U976 ( .A(\mem<27><6> ), .B(n1220), .Y(n1379) );
  OAI21X1 U977 ( .A(n102), .B(n1278), .C(n1379), .Y(n2274) );
  NAND2X1 U978 ( .A(\mem<27><7> ), .B(n1220), .Y(n1380) );
  OAI21X1 U979 ( .A(n102), .B(n1279), .C(n1380), .Y(n2273) );
  NAND2X1 U980 ( .A(\mem<27><8> ), .B(n1221), .Y(n1381) );
  OAI21X1 U981 ( .A(n102), .B(n1280), .C(n1381), .Y(n2272) );
  NAND2X1 U982 ( .A(\mem<27><9> ), .B(n1221), .Y(n1382) );
  OAI21X1 U983 ( .A(n102), .B(n1282), .C(n1382), .Y(n2271) );
  NAND2X1 U984 ( .A(\mem<27><10> ), .B(n1221), .Y(n1383) );
  OAI21X1 U985 ( .A(n102), .B(n1283), .C(n1383), .Y(n2270) );
  NAND2X1 U986 ( .A(\mem<27><11> ), .B(n1221), .Y(n1384) );
  OAI21X1 U987 ( .A(n102), .B(n1285), .C(n1384), .Y(n2269) );
  NAND2X1 U988 ( .A(\mem<27><12> ), .B(n1221), .Y(n1385) );
  OAI21X1 U989 ( .A(n102), .B(n1287), .C(n1385), .Y(n2268) );
  NAND2X1 U990 ( .A(\mem<27><13> ), .B(n1221), .Y(n1386) );
  OAI21X1 U991 ( .A(n102), .B(n1289), .C(n1386), .Y(n2267) );
  NAND2X1 U992 ( .A(\mem<27><14> ), .B(n1221), .Y(n1387) );
  OAI21X1 U993 ( .A(n102), .B(n1291), .C(n1387), .Y(n2266) );
  NAND2X1 U994 ( .A(\mem<27><15> ), .B(n1221), .Y(n1388) );
  OAI21X1 U995 ( .A(n102), .B(n1293), .C(n1388), .Y(n2265) );
  NAND3X1 U996 ( .A(n1299), .B(n1296), .C(n1295), .Y(n1389) );
  NAND2X1 U997 ( .A(\mem<26><0> ), .B(n1222), .Y(n1390) );
  OAI21X1 U998 ( .A(n104), .B(n1270), .C(n1390), .Y(n2264) );
  NAND2X1 U999 ( .A(\mem<26><1> ), .B(n1222), .Y(n1391) );
  OAI21X1 U1000 ( .A(n104), .B(n1272), .C(n1391), .Y(n2263) );
  NAND2X1 U1001 ( .A(\mem<26><2> ), .B(n1222), .Y(n1392) );
  OAI21X1 U1002 ( .A(n104), .B(n1273), .C(n1392), .Y(n2262) );
  NAND2X1 U1003 ( .A(\mem<26><3> ), .B(n1222), .Y(n1393) );
  OAI21X1 U1004 ( .A(n104), .B(n1274), .C(n1393), .Y(n2261) );
  NAND2X1 U1005 ( .A(\mem<26><4> ), .B(n1222), .Y(n1394) );
  OAI21X1 U1006 ( .A(n104), .B(n1275), .C(n1394), .Y(n2260) );
  NAND2X1 U1007 ( .A(\mem<26><5> ), .B(n1222), .Y(n1395) );
  OAI21X1 U1008 ( .A(n104), .B(n1277), .C(n1395), .Y(n2259) );
  NAND2X1 U1009 ( .A(\mem<26><6> ), .B(n1222), .Y(n1396) );
  OAI21X1 U1010 ( .A(n104), .B(n1278), .C(n1396), .Y(n2258) );
  NAND2X1 U1011 ( .A(\mem<26><7> ), .B(n1222), .Y(n1397) );
  OAI21X1 U1012 ( .A(n104), .B(n1279), .C(n1397), .Y(n2257) );
  NAND2X1 U1013 ( .A(\mem<26><8> ), .B(n1223), .Y(n1398) );
  OAI21X1 U1014 ( .A(n104), .B(n1280), .C(n1398), .Y(n2256) );
  NAND2X1 U1015 ( .A(\mem<26><9> ), .B(n1223), .Y(n1399) );
  OAI21X1 U1016 ( .A(n104), .B(n1281), .C(n1399), .Y(n2255) );
  NAND2X1 U1017 ( .A(\mem<26><10> ), .B(n1223), .Y(n1400) );
  OAI21X1 U1018 ( .A(n104), .B(n1283), .C(n1400), .Y(n2254) );
  NAND2X1 U1019 ( .A(\mem<26><11> ), .B(n1223), .Y(n1401) );
  OAI21X1 U1020 ( .A(n104), .B(n1284), .C(n1401), .Y(n2253) );
  NAND2X1 U1021 ( .A(\mem<26><12> ), .B(n1223), .Y(n1402) );
  OAI21X1 U1022 ( .A(n104), .B(n1286), .C(n1402), .Y(n2252) );
  NAND2X1 U1023 ( .A(\mem<26><13> ), .B(n1223), .Y(n1403) );
  OAI21X1 U1024 ( .A(n104), .B(n1288), .C(n1403), .Y(n2251) );
  NAND2X1 U1025 ( .A(\mem<26><14> ), .B(n1223), .Y(n1404) );
  OAI21X1 U1026 ( .A(n104), .B(n1290), .C(n1404), .Y(n2250) );
  NAND2X1 U1027 ( .A(\mem<26><15> ), .B(n1223), .Y(n1405) );
  OAI21X1 U1028 ( .A(n104), .B(n1292), .C(n1405), .Y(n2249) );
  NAND3X1 U1029 ( .A(N10), .B(n1299), .C(n1297), .Y(n1406) );
  NAND2X1 U1030 ( .A(\mem<25><0> ), .B(n1224), .Y(n1407) );
  OAI21X1 U1031 ( .A(n106), .B(n1270), .C(n1407), .Y(n2248) );
  NAND2X1 U1032 ( .A(\mem<25><1> ), .B(n1224), .Y(n1408) );
  OAI21X1 U1033 ( .A(n106), .B(n1271), .C(n1408), .Y(n2247) );
  NAND2X1 U1034 ( .A(\mem<25><2> ), .B(n1224), .Y(n1409) );
  OAI21X1 U1035 ( .A(n106), .B(n1273), .C(n1409), .Y(n2246) );
  NAND2X1 U1036 ( .A(\mem<25><3> ), .B(n1224), .Y(n1410) );
  OAI21X1 U1037 ( .A(n106), .B(n1274), .C(n1410), .Y(n2245) );
  NAND2X1 U1038 ( .A(\mem<25><4> ), .B(n1224), .Y(n1411) );
  OAI21X1 U1039 ( .A(n106), .B(n1275), .C(n1411), .Y(n2244) );
  NAND2X1 U1040 ( .A(\mem<25><5> ), .B(n1224), .Y(n1412) );
  OAI21X1 U1041 ( .A(n106), .B(n1276), .C(n1412), .Y(n2243) );
  NAND2X1 U1042 ( .A(\mem<25><6> ), .B(n1224), .Y(n1413) );
  OAI21X1 U1043 ( .A(n106), .B(n1278), .C(n1413), .Y(n2242) );
  NAND2X1 U1044 ( .A(\mem<25><7> ), .B(n1224), .Y(n1414) );
  OAI21X1 U1045 ( .A(n106), .B(n1279), .C(n1414), .Y(n2241) );
  NAND2X1 U1046 ( .A(\mem<25><8> ), .B(n1225), .Y(n1415) );
  OAI21X1 U1047 ( .A(n106), .B(n1280), .C(n1415), .Y(n2240) );
  NAND2X1 U1048 ( .A(\mem<25><9> ), .B(n1225), .Y(n1416) );
  OAI21X1 U1049 ( .A(n106), .B(n1282), .C(n1416), .Y(n2239) );
  NAND2X1 U1050 ( .A(\mem<25><10> ), .B(n1225), .Y(n1417) );
  OAI21X1 U1051 ( .A(n106), .B(n1283), .C(n1417), .Y(n2238) );
  NAND2X1 U1052 ( .A(\mem<25><11> ), .B(n1225), .Y(n1418) );
  OAI21X1 U1053 ( .A(n106), .B(n1285), .C(n1418), .Y(n2237) );
  NAND2X1 U1054 ( .A(\mem<25><12> ), .B(n1225), .Y(n1419) );
  OAI21X1 U1055 ( .A(n106), .B(n1287), .C(n1419), .Y(n2236) );
  NAND2X1 U1056 ( .A(\mem<25><13> ), .B(n1225), .Y(n1420) );
  OAI21X1 U1057 ( .A(n106), .B(n1289), .C(n1420), .Y(n2235) );
  NAND2X1 U1058 ( .A(\mem<25><14> ), .B(n1225), .Y(n1421) );
  OAI21X1 U1059 ( .A(n106), .B(n1291), .C(n1421), .Y(n2234) );
  NAND2X1 U1060 ( .A(\mem<25><15> ), .B(n1225), .Y(n1422) );
  OAI21X1 U1061 ( .A(n106), .B(n1293), .C(n1422), .Y(n2233) );
  NOR3X1 U1062 ( .A(N10), .B(n1296), .C(n1298), .Y(n1816) );
  NAND2X1 U1063 ( .A(\mem<24><0> ), .B(n1227), .Y(n1423) );
  OAI21X1 U1064 ( .A(n1226), .B(n1270), .C(n1423), .Y(n2232) );
  NAND2X1 U1065 ( .A(\mem<24><1> ), .B(n1227), .Y(n1424) );
  OAI21X1 U1066 ( .A(n1226), .B(n1271), .C(n1424), .Y(n2231) );
  NAND2X1 U1067 ( .A(\mem<24><2> ), .B(n1227), .Y(n1425) );
  OAI21X1 U1068 ( .A(n1226), .B(n1273), .C(n1425), .Y(n2230) );
  NAND2X1 U1069 ( .A(\mem<24><3> ), .B(n1227), .Y(n1426) );
  OAI21X1 U1070 ( .A(n1226), .B(n1274), .C(n1426), .Y(n2229) );
  NAND2X1 U1071 ( .A(\mem<24><4> ), .B(n1227), .Y(n1427) );
  OAI21X1 U1072 ( .A(n1226), .B(n1275), .C(n1427), .Y(n2228) );
  NAND2X1 U1073 ( .A(\mem<24><5> ), .B(n1227), .Y(n1428) );
  OAI21X1 U1074 ( .A(n1226), .B(n1276), .C(n1428), .Y(n2227) );
  NAND2X1 U1075 ( .A(\mem<24><6> ), .B(n1227), .Y(n1429) );
  OAI21X1 U1076 ( .A(n1226), .B(n1278), .C(n1429), .Y(n2226) );
  NAND2X1 U1077 ( .A(\mem<24><7> ), .B(n1227), .Y(n1430) );
  OAI21X1 U1078 ( .A(n1226), .B(n1279), .C(n1430), .Y(n2225) );
  NAND2X1 U1079 ( .A(\mem<24><8> ), .B(n1228), .Y(n1431) );
  OAI21X1 U1080 ( .A(n1226), .B(n1280), .C(n1431), .Y(n2224) );
  NAND2X1 U1081 ( .A(\mem<24><9> ), .B(n1228), .Y(n1432) );
  OAI21X1 U1082 ( .A(n1226), .B(n1281), .C(n1432), .Y(n2223) );
  NAND2X1 U1083 ( .A(\mem<24><10> ), .B(n1228), .Y(n1433) );
  OAI21X1 U1084 ( .A(n1226), .B(n1283), .C(n1433), .Y(n2222) );
  NAND2X1 U1085 ( .A(\mem<24><11> ), .B(n1228), .Y(n1434) );
  OAI21X1 U1086 ( .A(n1226), .B(n1284), .C(n1434), .Y(n2221) );
  NAND2X1 U1087 ( .A(\mem<24><12> ), .B(n1228), .Y(n1435) );
  OAI21X1 U1088 ( .A(n1226), .B(n1286), .C(n1435), .Y(n2220) );
  NAND2X1 U1089 ( .A(\mem<24><13> ), .B(n1228), .Y(n1436) );
  OAI21X1 U1090 ( .A(n1226), .B(n1288), .C(n1436), .Y(n2219) );
  NAND2X1 U1091 ( .A(\mem<24><14> ), .B(n1228), .Y(n1437) );
  OAI21X1 U1092 ( .A(n1226), .B(n1290), .C(n1437), .Y(n2218) );
  NAND2X1 U1093 ( .A(\mem<24><15> ), .B(n1228), .Y(n1438) );
  OAI21X1 U1094 ( .A(n1226), .B(n1292), .C(n1438), .Y(n2217) );
  NAND2X1 U1095 ( .A(\mem<23><0> ), .B(n1229), .Y(n1439) );
  OAI21X1 U1096 ( .A(n108), .B(n1270), .C(n1439), .Y(n2216) );
  NAND2X1 U1097 ( .A(\mem<23><1> ), .B(n1229), .Y(n1440) );
  OAI21X1 U1098 ( .A(n108), .B(n1272), .C(n1440), .Y(n2215) );
  NAND2X1 U1099 ( .A(\mem<23><2> ), .B(n1229), .Y(n1441) );
  OAI21X1 U1100 ( .A(n108), .B(n1273), .C(n1441), .Y(n2214) );
  NAND2X1 U1101 ( .A(\mem<23><3> ), .B(n1229), .Y(n1442) );
  OAI21X1 U1102 ( .A(n108), .B(n1274), .C(n1442), .Y(n2213) );
  NAND2X1 U1103 ( .A(\mem<23><4> ), .B(n1229), .Y(n1443) );
  OAI21X1 U1104 ( .A(n108), .B(n1275), .C(n1443), .Y(n2212) );
  NAND2X1 U1105 ( .A(\mem<23><5> ), .B(n1229), .Y(n1444) );
  OAI21X1 U1106 ( .A(n108), .B(n1277), .C(n1444), .Y(n2211) );
  NAND2X1 U1107 ( .A(\mem<23><6> ), .B(n1229), .Y(n1445) );
  OAI21X1 U1108 ( .A(n108), .B(n1278), .C(n1445), .Y(n2210) );
  NAND2X1 U1109 ( .A(\mem<23><7> ), .B(n1229), .Y(n1446) );
  OAI21X1 U1110 ( .A(n108), .B(n1279), .C(n1446), .Y(n2209) );
  NAND2X1 U1111 ( .A(\mem<23><8> ), .B(n1230), .Y(n1447) );
  OAI21X1 U1112 ( .A(n108), .B(n1280), .C(n1447), .Y(n2208) );
  NAND2X1 U1113 ( .A(\mem<23><9> ), .B(n1230), .Y(n1448) );
  OAI21X1 U1114 ( .A(n108), .B(n1282), .C(n1448), .Y(n2207) );
  NAND2X1 U1115 ( .A(\mem<23><10> ), .B(n1230), .Y(n1449) );
  OAI21X1 U1116 ( .A(n108), .B(n1283), .C(n1449), .Y(n2206) );
  NAND2X1 U1117 ( .A(\mem<23><11> ), .B(n1230), .Y(n1450) );
  OAI21X1 U1118 ( .A(n108), .B(n1285), .C(n1450), .Y(n2205) );
  NAND2X1 U1119 ( .A(\mem<23><12> ), .B(n1230), .Y(n1451) );
  OAI21X1 U1120 ( .A(n108), .B(n1287), .C(n1451), .Y(n2204) );
  NAND2X1 U1121 ( .A(\mem<23><13> ), .B(n1230), .Y(n1452) );
  OAI21X1 U1122 ( .A(n108), .B(n1289), .C(n1452), .Y(n2203) );
  NAND2X1 U1123 ( .A(\mem<23><14> ), .B(n1230), .Y(n1453) );
  OAI21X1 U1124 ( .A(n108), .B(n1291), .C(n1453), .Y(n2202) );
  NAND2X1 U1125 ( .A(\mem<23><15> ), .B(n1230), .Y(n1454) );
  OAI21X1 U1126 ( .A(n108), .B(n1293), .C(n1454), .Y(n2201) );
  NAND2X1 U1127 ( .A(\mem<22><0> ), .B(n1231), .Y(n1455) );
  OAI21X1 U1128 ( .A(n110), .B(n1270), .C(n1455), .Y(n2200) );
  NAND2X1 U1129 ( .A(\mem<22><1> ), .B(n1231), .Y(n1456) );
  OAI21X1 U1130 ( .A(n110), .B(n1272), .C(n1456), .Y(n2199) );
  NAND2X1 U1131 ( .A(\mem<22><2> ), .B(n1231), .Y(n1457) );
  OAI21X1 U1132 ( .A(n110), .B(n1273), .C(n1457), .Y(n2198) );
  NAND2X1 U1133 ( .A(\mem<22><3> ), .B(n1231), .Y(n1458) );
  OAI21X1 U1134 ( .A(n110), .B(n1274), .C(n1458), .Y(n2197) );
  NAND2X1 U1135 ( .A(\mem<22><4> ), .B(n1231), .Y(n1459) );
  OAI21X1 U1136 ( .A(n110), .B(n1275), .C(n1459), .Y(n2196) );
  NAND2X1 U1137 ( .A(\mem<22><5> ), .B(n1231), .Y(n1460) );
  OAI21X1 U1138 ( .A(n110), .B(n1277), .C(n1460), .Y(n2195) );
  NAND2X1 U1139 ( .A(\mem<22><6> ), .B(n1231), .Y(n1461) );
  OAI21X1 U1140 ( .A(n110), .B(n1278), .C(n1461), .Y(n2194) );
  NAND2X1 U1141 ( .A(\mem<22><7> ), .B(n1231), .Y(n1462) );
  OAI21X1 U1142 ( .A(n110), .B(n1279), .C(n1462), .Y(n2193) );
  NAND2X1 U1143 ( .A(\mem<22><8> ), .B(n1232), .Y(n1463) );
  OAI21X1 U1144 ( .A(n110), .B(n1280), .C(n1463), .Y(n2192) );
  NAND2X1 U1145 ( .A(\mem<22><9> ), .B(n1232), .Y(n1464) );
  OAI21X1 U1146 ( .A(n110), .B(n1282), .C(n1464), .Y(n2191) );
  NAND2X1 U1147 ( .A(\mem<22><10> ), .B(n1232), .Y(n1465) );
  OAI21X1 U1148 ( .A(n110), .B(n1283), .C(n1465), .Y(n2190) );
  NAND2X1 U1149 ( .A(\mem<22><11> ), .B(n1232), .Y(n1466) );
  OAI21X1 U1150 ( .A(n110), .B(n1285), .C(n1466), .Y(n2189) );
  NAND2X1 U1151 ( .A(\mem<22><12> ), .B(n1232), .Y(n1467) );
  OAI21X1 U1152 ( .A(n110), .B(n1287), .C(n1467), .Y(n2188) );
  NAND2X1 U1153 ( .A(\mem<22><13> ), .B(n1232), .Y(n1468) );
  OAI21X1 U1154 ( .A(n110), .B(n1289), .C(n1468), .Y(n2187) );
  NAND2X1 U1155 ( .A(\mem<22><14> ), .B(n1232), .Y(n1469) );
  OAI21X1 U1156 ( .A(n110), .B(n1291), .C(n1469), .Y(n2186) );
  NAND2X1 U1157 ( .A(\mem<22><15> ), .B(n1232), .Y(n1470) );
  OAI21X1 U1158 ( .A(n110), .B(n1293), .C(n1470), .Y(n2185) );
  NAND2X1 U1159 ( .A(\mem<21><0> ), .B(n1233), .Y(n1471) );
  OAI21X1 U1160 ( .A(n112), .B(n1270), .C(n1471), .Y(n2184) );
  NAND2X1 U1161 ( .A(\mem<21><1> ), .B(n1233), .Y(n1472) );
  OAI21X1 U1162 ( .A(n112), .B(n1272), .C(n1472), .Y(n2183) );
  NAND2X1 U1163 ( .A(\mem<21><2> ), .B(n1233), .Y(n1473) );
  OAI21X1 U1164 ( .A(n112), .B(n1273), .C(n1473), .Y(n2182) );
  NAND2X1 U1165 ( .A(\mem<21><3> ), .B(n1233), .Y(n1474) );
  OAI21X1 U1166 ( .A(n112), .B(n1274), .C(n1474), .Y(n2181) );
  NAND2X1 U1167 ( .A(\mem<21><4> ), .B(n1233), .Y(n1475) );
  OAI21X1 U1168 ( .A(n112), .B(n1275), .C(n1475), .Y(n2180) );
  NAND2X1 U1169 ( .A(\mem<21><5> ), .B(n1233), .Y(n1476) );
  OAI21X1 U1170 ( .A(n112), .B(n1277), .C(n1476), .Y(n2179) );
  NAND2X1 U1171 ( .A(\mem<21><6> ), .B(n1233), .Y(n1477) );
  OAI21X1 U1172 ( .A(n112), .B(n1278), .C(n1477), .Y(n2178) );
  NAND2X1 U1173 ( .A(\mem<21><7> ), .B(n1233), .Y(n1478) );
  OAI21X1 U1174 ( .A(n112), .B(n1279), .C(n1478), .Y(n2177) );
  NAND2X1 U1175 ( .A(\mem<21><8> ), .B(n1234), .Y(n1479) );
  OAI21X1 U1177 ( .A(n112), .B(n1280), .C(n1479), .Y(n2176) );
  NAND2X1 U1178 ( .A(\mem<21><9> ), .B(n1234), .Y(n1480) );
  OAI21X1 U1179 ( .A(n112), .B(n1282), .C(n1480), .Y(n2175) );
  NAND2X1 U1180 ( .A(\mem<21><10> ), .B(n1234), .Y(n1481) );
  OAI21X1 U1181 ( .A(n112), .B(n1283), .C(n1481), .Y(n2174) );
  NAND2X1 U1182 ( .A(\mem<21><11> ), .B(n1234), .Y(n1482) );
  OAI21X1 U1183 ( .A(n112), .B(n1285), .C(n1482), .Y(n2173) );
  NAND2X1 U1184 ( .A(\mem<21><12> ), .B(n1234), .Y(n1483) );
  OAI21X1 U1185 ( .A(n112), .B(n1287), .C(n1483), .Y(n2172) );
  NAND2X1 U1186 ( .A(\mem<21><13> ), .B(n1234), .Y(n1484) );
  OAI21X1 U1187 ( .A(n112), .B(n1289), .C(n1484), .Y(n2171) );
  NAND2X1 U1188 ( .A(\mem<21><14> ), .B(n1234), .Y(n1485) );
  OAI21X1 U1189 ( .A(n112), .B(n1291), .C(n1485), .Y(n2170) );
  NAND2X1 U1190 ( .A(\mem<21><15> ), .B(n1234), .Y(n1486) );
  OAI21X1 U1191 ( .A(n112), .B(n1293), .C(n1486), .Y(n2169) );
  NAND2X1 U1192 ( .A(\mem<20><0> ), .B(n1235), .Y(n1487) );
  OAI21X1 U1193 ( .A(n114), .B(n1270), .C(n1487), .Y(n2168) );
  NAND2X1 U1194 ( .A(\mem<20><1> ), .B(n1235), .Y(n1488) );
  OAI21X1 U1195 ( .A(n114), .B(n1272), .C(n1488), .Y(n2167) );
  NAND2X1 U1196 ( .A(\mem<20><2> ), .B(n1235), .Y(n1489) );
  OAI21X1 U1197 ( .A(n114), .B(n1273), .C(n1489), .Y(n2166) );
  NAND2X1 U1198 ( .A(\mem<20><3> ), .B(n1235), .Y(n1490) );
  OAI21X1 U1199 ( .A(n114), .B(n1274), .C(n1490), .Y(n2165) );
  NAND2X1 U1200 ( .A(\mem<20><4> ), .B(n1235), .Y(n1491) );
  OAI21X1 U1201 ( .A(n114), .B(n1275), .C(n1491), .Y(n2164) );
  NAND2X1 U1202 ( .A(\mem<20><5> ), .B(n1235), .Y(n1492) );
  OAI21X1 U1203 ( .A(n114), .B(n1277), .C(n1492), .Y(n2163) );
  NAND2X1 U1204 ( .A(\mem<20><6> ), .B(n1235), .Y(n1493) );
  OAI21X1 U1205 ( .A(n114), .B(n1278), .C(n1493), .Y(n2162) );
  NAND2X1 U1206 ( .A(\mem<20><7> ), .B(n1235), .Y(n1494) );
  OAI21X1 U1207 ( .A(n114), .B(n1279), .C(n1494), .Y(n2161) );
  NAND2X1 U1208 ( .A(\mem<20><8> ), .B(n1236), .Y(n1495) );
  OAI21X1 U1209 ( .A(n114), .B(n1280), .C(n1495), .Y(n2160) );
  NAND2X1 U1210 ( .A(\mem<20><9> ), .B(n1236), .Y(n1496) );
  OAI21X1 U1211 ( .A(n114), .B(n1282), .C(n1496), .Y(n2159) );
  NAND2X1 U1212 ( .A(\mem<20><10> ), .B(n1236), .Y(n1497) );
  OAI21X1 U1213 ( .A(n114), .B(n1283), .C(n1497), .Y(n2158) );
  NAND2X1 U1214 ( .A(\mem<20><11> ), .B(n1236), .Y(n1498) );
  OAI21X1 U1215 ( .A(n114), .B(n1285), .C(n1498), .Y(n2157) );
  NAND2X1 U1216 ( .A(\mem<20><12> ), .B(n1236), .Y(n1499) );
  OAI21X1 U1217 ( .A(n114), .B(n1287), .C(n1499), .Y(n2156) );
  NAND2X1 U1218 ( .A(\mem<20><13> ), .B(n1236), .Y(n1500) );
  OAI21X1 U1219 ( .A(n114), .B(n1289), .C(n1500), .Y(n2155) );
  NAND2X1 U1220 ( .A(\mem<20><14> ), .B(n1236), .Y(n1501) );
  OAI21X1 U1221 ( .A(n114), .B(n1291), .C(n1501), .Y(n2154) );
  NAND2X1 U1222 ( .A(\mem<20><15> ), .B(n1236), .Y(n1502) );
  OAI21X1 U1223 ( .A(n114), .B(n1293), .C(n1502), .Y(n2153) );
  NAND2X1 U1224 ( .A(\mem<19><0> ), .B(n1237), .Y(n1503) );
  OAI21X1 U1225 ( .A(n116), .B(n1270), .C(n1503), .Y(n2152) );
  NAND2X1 U1226 ( .A(\mem<19><1> ), .B(n1237), .Y(n1504) );
  OAI21X1 U1227 ( .A(n116), .B(n1272), .C(n1504), .Y(n2151) );
  NAND2X1 U1228 ( .A(\mem<19><2> ), .B(n1237), .Y(n1505) );
  OAI21X1 U1229 ( .A(n116), .B(n1273), .C(n1505), .Y(n2150) );
  NAND2X1 U1230 ( .A(\mem<19><3> ), .B(n1237), .Y(n1506) );
  OAI21X1 U1231 ( .A(n116), .B(n1274), .C(n1506), .Y(n2149) );
  NAND2X1 U1232 ( .A(\mem<19><4> ), .B(n1237), .Y(n1507) );
  OAI21X1 U1233 ( .A(n116), .B(n1275), .C(n1507), .Y(n2148) );
  NAND2X1 U1234 ( .A(\mem<19><5> ), .B(n1237), .Y(n1508) );
  OAI21X1 U1235 ( .A(n116), .B(n1277), .C(n1508), .Y(n2147) );
  NAND2X1 U1236 ( .A(\mem<19><6> ), .B(n1237), .Y(n1509) );
  OAI21X1 U1237 ( .A(n116), .B(n1278), .C(n1509), .Y(n2146) );
  NAND2X1 U1238 ( .A(\mem<19><7> ), .B(n1237), .Y(n1510) );
  OAI21X1 U1239 ( .A(n116), .B(n1279), .C(n1510), .Y(n2145) );
  NAND2X1 U1240 ( .A(\mem<19><8> ), .B(n1238), .Y(n1511) );
  OAI21X1 U1241 ( .A(n116), .B(n1280), .C(n1511), .Y(n2144) );
  NAND2X1 U1242 ( .A(\mem<19><9> ), .B(n1238), .Y(n1512) );
  OAI21X1 U1243 ( .A(n116), .B(n1282), .C(n1512), .Y(n2143) );
  NAND2X1 U1244 ( .A(\mem<19><10> ), .B(n1238), .Y(n1513) );
  OAI21X1 U1245 ( .A(n116), .B(n1283), .C(n1513), .Y(n2142) );
  NAND2X1 U1246 ( .A(\mem<19><11> ), .B(n1238), .Y(n1514) );
  OAI21X1 U1247 ( .A(n116), .B(n1285), .C(n1514), .Y(n2141) );
  NAND2X1 U1248 ( .A(\mem<19><12> ), .B(n1238), .Y(n1515) );
  OAI21X1 U1249 ( .A(n116), .B(n1287), .C(n1515), .Y(n2140) );
  NAND2X1 U1250 ( .A(\mem<19><13> ), .B(n1238), .Y(n1516) );
  OAI21X1 U1251 ( .A(n116), .B(n1289), .C(n1516), .Y(n2139) );
  NAND2X1 U1252 ( .A(\mem<19><14> ), .B(n1238), .Y(n1517) );
  OAI21X1 U1253 ( .A(n116), .B(n1291), .C(n1517), .Y(n2138) );
  NAND2X1 U1254 ( .A(\mem<19><15> ), .B(n1238), .Y(n1518) );
  OAI21X1 U1255 ( .A(n116), .B(n1293), .C(n1518), .Y(n2137) );
  NAND2X1 U1256 ( .A(\mem<18><0> ), .B(n1239), .Y(n1519) );
  OAI21X1 U1257 ( .A(n118), .B(n1270), .C(n1519), .Y(n2136) );
  NAND2X1 U1258 ( .A(\mem<18><1> ), .B(n1239), .Y(n1520) );
  OAI21X1 U1259 ( .A(n118), .B(n1272), .C(n1520), .Y(n2135) );
  NAND2X1 U1260 ( .A(\mem<18><2> ), .B(n1239), .Y(n1521) );
  OAI21X1 U1261 ( .A(n118), .B(n1273), .C(n1521), .Y(n2134) );
  NAND2X1 U1262 ( .A(\mem<18><3> ), .B(n1239), .Y(n1522) );
  OAI21X1 U1263 ( .A(n118), .B(n1274), .C(n1522), .Y(n2133) );
  NAND2X1 U1264 ( .A(\mem<18><4> ), .B(n1239), .Y(n1523) );
  OAI21X1 U1265 ( .A(n118), .B(n1275), .C(n1523), .Y(n2132) );
  NAND2X1 U1266 ( .A(\mem<18><5> ), .B(n1239), .Y(n1524) );
  OAI21X1 U1267 ( .A(n118), .B(n1277), .C(n1524), .Y(n2131) );
  NAND2X1 U1268 ( .A(\mem<18><6> ), .B(n1239), .Y(n1525) );
  OAI21X1 U1269 ( .A(n118), .B(n1278), .C(n1525), .Y(n2130) );
  NAND2X1 U1270 ( .A(\mem<18><7> ), .B(n1239), .Y(n1526) );
  OAI21X1 U1271 ( .A(n118), .B(n1279), .C(n1526), .Y(n2129) );
  NAND2X1 U1272 ( .A(\mem<18><8> ), .B(n1240), .Y(n1527) );
  OAI21X1 U1273 ( .A(n118), .B(n1280), .C(n1527), .Y(n2128) );
  NAND2X1 U1274 ( .A(\mem<18><9> ), .B(n1240), .Y(n1528) );
  OAI21X1 U1275 ( .A(n118), .B(n1282), .C(n1528), .Y(n2127) );
  NAND2X1 U1276 ( .A(\mem<18><10> ), .B(n1240), .Y(n1529) );
  OAI21X1 U1277 ( .A(n118), .B(n1283), .C(n1529), .Y(n2126) );
  NAND2X1 U1278 ( .A(\mem<18><11> ), .B(n1240), .Y(n1530) );
  OAI21X1 U1279 ( .A(n118), .B(n1285), .C(n1530), .Y(n2125) );
  NAND2X1 U1280 ( .A(\mem<18><12> ), .B(n1240), .Y(n1531) );
  OAI21X1 U1281 ( .A(n118), .B(n1287), .C(n1531), .Y(n2124) );
  NAND2X1 U1282 ( .A(\mem<18><13> ), .B(n1240), .Y(n1532) );
  OAI21X1 U1283 ( .A(n118), .B(n1289), .C(n1532), .Y(n2123) );
  NAND2X1 U1284 ( .A(\mem<18><14> ), .B(n1240), .Y(n1533) );
  OAI21X1 U1285 ( .A(n118), .B(n1291), .C(n1533), .Y(n2122) );
  NAND2X1 U1286 ( .A(\mem<18><15> ), .B(n1240), .Y(n1534) );
  OAI21X1 U1287 ( .A(n118), .B(n1293), .C(n1534), .Y(n2121) );
  NAND2X1 U1288 ( .A(\mem<17><0> ), .B(n1241), .Y(n1535) );
  OAI21X1 U1289 ( .A(n120), .B(n1270), .C(n1535), .Y(n2120) );
  NAND2X1 U1290 ( .A(\mem<17><1> ), .B(n1241), .Y(n1536) );
  OAI21X1 U1291 ( .A(n120), .B(n1272), .C(n1536), .Y(n2119) );
  NAND2X1 U1292 ( .A(\mem<17><2> ), .B(n1241), .Y(n1537) );
  OAI21X1 U1293 ( .A(n120), .B(n1273), .C(n1537), .Y(n2118) );
  NAND2X1 U1294 ( .A(\mem<17><3> ), .B(n1241), .Y(n1538) );
  OAI21X1 U1295 ( .A(n120), .B(n1274), .C(n1538), .Y(n2117) );
  NAND2X1 U1296 ( .A(\mem<17><4> ), .B(n1241), .Y(n1539) );
  OAI21X1 U1297 ( .A(n120), .B(n1275), .C(n1539), .Y(n2116) );
  NAND2X1 U1298 ( .A(\mem<17><5> ), .B(n1241), .Y(n1540) );
  OAI21X1 U1299 ( .A(n120), .B(n1277), .C(n1540), .Y(n2115) );
  NAND2X1 U1300 ( .A(\mem<17><6> ), .B(n1241), .Y(n1541) );
  OAI21X1 U1301 ( .A(n120), .B(n1278), .C(n1541), .Y(n2114) );
  NAND2X1 U1302 ( .A(\mem<17><7> ), .B(n1241), .Y(n1542) );
  OAI21X1 U1303 ( .A(n120), .B(n1279), .C(n1542), .Y(n2113) );
  NAND2X1 U1304 ( .A(\mem<17><8> ), .B(n1242), .Y(n1543) );
  OAI21X1 U1305 ( .A(n120), .B(n1280), .C(n1543), .Y(n2112) );
  NAND2X1 U1306 ( .A(\mem<17><9> ), .B(n1242), .Y(n1544) );
  OAI21X1 U1307 ( .A(n120), .B(n1282), .C(n1544), .Y(n2111) );
  NAND2X1 U1308 ( .A(\mem<17><10> ), .B(n1242), .Y(n1545) );
  OAI21X1 U1309 ( .A(n120), .B(n1283), .C(n1545), .Y(n2110) );
  NAND2X1 U1310 ( .A(\mem<17><11> ), .B(n1242), .Y(n1546) );
  OAI21X1 U1311 ( .A(n120), .B(n1285), .C(n1546), .Y(n2109) );
  NAND2X1 U1312 ( .A(\mem<17><12> ), .B(n1242), .Y(n1547) );
  OAI21X1 U1313 ( .A(n120), .B(n1287), .C(n1547), .Y(n2108) );
  NAND2X1 U1314 ( .A(\mem<17><13> ), .B(n1242), .Y(n1548) );
  OAI21X1 U1315 ( .A(n120), .B(n1289), .C(n1548), .Y(n2107) );
  NAND2X1 U1316 ( .A(\mem<17><14> ), .B(n1242), .Y(n1549) );
  OAI21X1 U1317 ( .A(n120), .B(n1291), .C(n1549), .Y(n2106) );
  NAND2X1 U1318 ( .A(\mem<17><15> ), .B(n1242), .Y(n1550) );
  OAI21X1 U1319 ( .A(n120), .B(n1293), .C(n1550), .Y(n2105) );
  NAND2X1 U1320 ( .A(\mem<16><0> ), .B(n1244), .Y(n1551) );
  OAI21X1 U1321 ( .A(n1243), .B(n1270), .C(n1551), .Y(n2104) );
  NAND2X1 U1322 ( .A(\mem<16><1> ), .B(n1244), .Y(n1552) );
  OAI21X1 U1323 ( .A(n1243), .B(n1272), .C(n1552), .Y(n2103) );
  NAND2X1 U1324 ( .A(\mem<16><2> ), .B(n1244), .Y(n1553) );
  OAI21X1 U1325 ( .A(n1243), .B(n1273), .C(n1553), .Y(n2102) );
  NAND2X1 U1326 ( .A(\mem<16><3> ), .B(n1244), .Y(n1554) );
  OAI21X1 U1327 ( .A(n1243), .B(n1274), .C(n1554), .Y(n2101) );
  NAND2X1 U1328 ( .A(\mem<16><4> ), .B(n1244), .Y(n1555) );
  OAI21X1 U1329 ( .A(n1243), .B(n1275), .C(n1555), .Y(n2100) );
  NAND2X1 U1330 ( .A(\mem<16><5> ), .B(n1244), .Y(n1556) );
  OAI21X1 U1331 ( .A(n1243), .B(n1277), .C(n1556), .Y(n2099) );
  NAND2X1 U1332 ( .A(\mem<16><6> ), .B(n1244), .Y(n1557) );
  OAI21X1 U1333 ( .A(n1243), .B(n1278), .C(n1557), .Y(n2098) );
  NAND2X1 U1334 ( .A(\mem<16><7> ), .B(n1244), .Y(n1558) );
  OAI21X1 U1335 ( .A(n1243), .B(n1279), .C(n1558), .Y(n2097) );
  NAND2X1 U1336 ( .A(\mem<16><8> ), .B(n1245), .Y(n1559) );
  OAI21X1 U1337 ( .A(n1243), .B(n1280), .C(n1559), .Y(n2096) );
  NAND2X1 U1338 ( .A(\mem<16><9> ), .B(n1245), .Y(n1560) );
  OAI21X1 U1339 ( .A(n1243), .B(n1282), .C(n1560), .Y(n2095) );
  NAND2X1 U1340 ( .A(\mem<16><10> ), .B(n1245), .Y(n1561) );
  OAI21X1 U1341 ( .A(n1243), .B(n1283), .C(n1561), .Y(n2094) );
  NAND2X1 U1342 ( .A(\mem<16><11> ), .B(n1245), .Y(n1562) );
  OAI21X1 U1343 ( .A(n1243), .B(n1285), .C(n1562), .Y(n2093) );
  NAND2X1 U1344 ( .A(\mem<16><12> ), .B(n1245), .Y(n1563) );
  OAI21X1 U1345 ( .A(n1243), .B(n1287), .C(n1563), .Y(n2092) );
  NAND2X1 U1346 ( .A(\mem<16><13> ), .B(n1245), .Y(n1564) );
  OAI21X1 U1347 ( .A(n1243), .B(n1289), .C(n1564), .Y(n2091) );
  NAND2X1 U1348 ( .A(\mem<16><14> ), .B(n1245), .Y(n1565) );
  OAI21X1 U1349 ( .A(n1243), .B(n1291), .C(n1565), .Y(n2090) );
  NAND2X1 U1350 ( .A(\mem<16><15> ), .B(n1245), .Y(n1566) );
  OAI21X1 U1351 ( .A(n1243), .B(n1293), .C(n1566), .Y(n2089) );
  NAND3X1 U1352 ( .A(n1300), .B(n2345), .C(n1303), .Y(n1567) );
  NAND2X1 U1353 ( .A(\mem<15><0> ), .B(n1246), .Y(n1568) );
  OAI21X1 U1354 ( .A(n122), .B(n1270), .C(n1568), .Y(n2088) );
  NAND2X1 U1355 ( .A(\mem<15><1> ), .B(n1246), .Y(n1569) );
  OAI21X1 U1356 ( .A(n122), .B(n1272), .C(n1569), .Y(n2087) );
  NAND2X1 U1357 ( .A(\mem<15><2> ), .B(n1246), .Y(n1570) );
  OAI21X1 U1358 ( .A(n122), .B(n1273), .C(n1570), .Y(n2086) );
  NAND2X1 U1359 ( .A(\mem<15><3> ), .B(n1246), .Y(n1571) );
  OAI21X1 U1360 ( .A(n122), .B(n1274), .C(n1571), .Y(n2085) );
  NAND2X1 U1361 ( .A(\mem<15><4> ), .B(n1246), .Y(n1572) );
  OAI21X1 U1362 ( .A(n122), .B(n1275), .C(n1572), .Y(n2084) );
  NAND2X1 U1363 ( .A(\mem<15><5> ), .B(n1246), .Y(n1573) );
  OAI21X1 U1364 ( .A(n122), .B(n1277), .C(n1573), .Y(n2083) );
  NAND2X1 U1365 ( .A(\mem<15><6> ), .B(n1246), .Y(n1574) );
  OAI21X1 U1366 ( .A(n122), .B(n1278), .C(n1574), .Y(n2082) );
  NAND2X1 U1367 ( .A(\mem<15><7> ), .B(n1246), .Y(n1575) );
  OAI21X1 U1368 ( .A(n122), .B(n1279), .C(n1575), .Y(n2081) );
  NAND2X1 U1369 ( .A(\mem<15><8> ), .B(n1247), .Y(n1576) );
  OAI21X1 U1370 ( .A(n122), .B(n1280), .C(n1576), .Y(n2080) );
  NAND2X1 U1371 ( .A(\mem<15><9> ), .B(n1247), .Y(n1577) );
  OAI21X1 U1372 ( .A(n122), .B(n1282), .C(n1577), .Y(n2079) );
  NAND2X1 U1373 ( .A(\mem<15><10> ), .B(n1247), .Y(n1578) );
  OAI21X1 U1374 ( .A(n122), .B(n1283), .C(n1578), .Y(n2078) );
  NAND2X1 U1375 ( .A(\mem<15><11> ), .B(n1247), .Y(n1579) );
  OAI21X1 U1376 ( .A(n122), .B(n1285), .C(n1579), .Y(n2077) );
  NAND2X1 U1377 ( .A(\mem<15><12> ), .B(n1247), .Y(n1580) );
  OAI21X1 U1378 ( .A(n122), .B(n1287), .C(n1580), .Y(n2076) );
  NAND2X1 U1379 ( .A(\mem<15><13> ), .B(n1247), .Y(n1581) );
  OAI21X1 U1380 ( .A(n122), .B(n1289), .C(n1581), .Y(n2075) );
  NAND2X1 U1381 ( .A(\mem<15><14> ), .B(n1247), .Y(n1582) );
  OAI21X1 U1382 ( .A(n122), .B(n1291), .C(n1582), .Y(n2074) );
  NAND2X1 U1383 ( .A(\mem<15><15> ), .B(n1247), .Y(n1583) );
  OAI21X1 U1384 ( .A(n122), .B(n1293), .C(n1583), .Y(n2073) );
  NAND2X1 U1385 ( .A(\mem<14><0> ), .B(n1248), .Y(n1584) );
  OAI21X1 U1386 ( .A(n124), .B(n1270), .C(n1584), .Y(n2072) );
  NAND2X1 U1387 ( .A(\mem<14><1> ), .B(n1248), .Y(n1585) );
  OAI21X1 U1388 ( .A(n124), .B(n1272), .C(n1585), .Y(n2071) );
  NAND2X1 U1389 ( .A(\mem<14><2> ), .B(n1248), .Y(n1586) );
  OAI21X1 U1390 ( .A(n124), .B(n1273), .C(n1586), .Y(n2070) );
  NAND2X1 U1391 ( .A(\mem<14><3> ), .B(n1248), .Y(n1587) );
  OAI21X1 U1392 ( .A(n124), .B(n1274), .C(n1587), .Y(n2069) );
  NAND2X1 U1393 ( .A(\mem<14><4> ), .B(n1248), .Y(n1588) );
  OAI21X1 U1394 ( .A(n124), .B(n1275), .C(n1588), .Y(n2068) );
  NAND2X1 U1395 ( .A(\mem<14><5> ), .B(n1248), .Y(n1589) );
  OAI21X1 U1396 ( .A(n124), .B(n1277), .C(n1589), .Y(n2067) );
  NAND2X1 U1397 ( .A(\mem<14><6> ), .B(n1248), .Y(n1590) );
  OAI21X1 U1398 ( .A(n124), .B(n1278), .C(n1590), .Y(n2066) );
  NAND2X1 U1399 ( .A(\mem<14><7> ), .B(n1248), .Y(n1591) );
  OAI21X1 U1400 ( .A(n124), .B(n1279), .C(n1591), .Y(n2065) );
  NAND2X1 U1401 ( .A(\mem<14><8> ), .B(n1249), .Y(n1592) );
  OAI21X1 U1402 ( .A(n124), .B(n1280), .C(n1592), .Y(n2064) );
  NAND2X1 U1403 ( .A(\mem<14><9> ), .B(n1249), .Y(n1593) );
  OAI21X1 U1404 ( .A(n124), .B(n1282), .C(n1593), .Y(n2063) );
  NAND2X1 U1405 ( .A(\mem<14><10> ), .B(n1249), .Y(n1594) );
  OAI21X1 U1406 ( .A(n124), .B(n1283), .C(n1594), .Y(n2062) );
  NAND2X1 U1407 ( .A(\mem<14><11> ), .B(n1249), .Y(n1595) );
  OAI21X1 U1408 ( .A(n124), .B(n1285), .C(n1595), .Y(n2061) );
  NAND2X1 U1409 ( .A(\mem<14><12> ), .B(n1249), .Y(n1596) );
  OAI21X1 U1410 ( .A(n124), .B(n1287), .C(n1596), .Y(n2060) );
  NAND2X1 U1411 ( .A(\mem<14><13> ), .B(n1249), .Y(n1597) );
  OAI21X1 U1412 ( .A(n124), .B(n1289), .C(n1597), .Y(n2059) );
  NAND2X1 U1413 ( .A(\mem<14><14> ), .B(n1249), .Y(n1598) );
  OAI21X1 U1414 ( .A(n124), .B(n1291), .C(n1598), .Y(n2058) );
  NAND2X1 U1415 ( .A(\mem<14><15> ), .B(n1249), .Y(n1599) );
  OAI21X1 U1416 ( .A(n124), .B(n1293), .C(n1599), .Y(n2057) );
  NAND2X1 U1417 ( .A(\mem<13><0> ), .B(n1250), .Y(n1600) );
  OAI21X1 U1418 ( .A(n126), .B(n1270), .C(n1600), .Y(n2056) );
  NAND2X1 U1419 ( .A(\mem<13><1> ), .B(n1250), .Y(n1601) );
  OAI21X1 U1420 ( .A(n126), .B(n1272), .C(n1601), .Y(n2055) );
  NAND2X1 U1421 ( .A(\mem<13><2> ), .B(n1250), .Y(n1602) );
  OAI21X1 U1422 ( .A(n126), .B(n1273), .C(n1602), .Y(n2054) );
  NAND2X1 U1423 ( .A(\mem<13><3> ), .B(n1250), .Y(n1603) );
  OAI21X1 U1424 ( .A(n126), .B(n1274), .C(n1603), .Y(n2053) );
  NAND2X1 U1425 ( .A(\mem<13><4> ), .B(n1250), .Y(n1604) );
  OAI21X1 U1426 ( .A(n126), .B(n1275), .C(n1604), .Y(n2052) );
  NAND2X1 U1427 ( .A(\mem<13><5> ), .B(n1250), .Y(n1605) );
  OAI21X1 U1428 ( .A(n126), .B(n1277), .C(n1605), .Y(n2051) );
  NAND2X1 U1429 ( .A(\mem<13><6> ), .B(n1250), .Y(n1606) );
  OAI21X1 U1430 ( .A(n126), .B(n1278), .C(n1606), .Y(n2050) );
  NAND2X1 U1431 ( .A(\mem<13><7> ), .B(n1250), .Y(n1607) );
  OAI21X1 U1432 ( .A(n126), .B(n1279), .C(n1607), .Y(n2049) );
  NAND2X1 U1433 ( .A(\mem<13><8> ), .B(n1251), .Y(n1608) );
  OAI21X1 U1434 ( .A(n126), .B(n1280), .C(n1608), .Y(n2048) );
  NAND2X1 U1435 ( .A(\mem<13><9> ), .B(n1251), .Y(n1609) );
  OAI21X1 U1436 ( .A(n126), .B(n1282), .C(n1609), .Y(n2047) );
  NAND2X1 U1437 ( .A(\mem<13><10> ), .B(n1251), .Y(n1610) );
  OAI21X1 U1438 ( .A(n126), .B(n1283), .C(n1610), .Y(n2046) );
  NAND2X1 U1439 ( .A(\mem<13><11> ), .B(n1251), .Y(n1611) );
  OAI21X1 U1440 ( .A(n126), .B(n1285), .C(n1611), .Y(n2045) );
  NAND2X1 U1441 ( .A(\mem<13><12> ), .B(n1251), .Y(n1612) );
  OAI21X1 U1442 ( .A(n126), .B(n1287), .C(n1612), .Y(n2044) );
  NAND2X1 U1443 ( .A(\mem<13><13> ), .B(n1251), .Y(n1613) );
  OAI21X1 U1444 ( .A(n126), .B(n1289), .C(n1613), .Y(n2043) );
  NAND2X1 U1445 ( .A(\mem<13><14> ), .B(n1251), .Y(n1614) );
  OAI21X1 U1446 ( .A(n126), .B(n1291), .C(n1614), .Y(n2042) );
  NAND2X1 U1447 ( .A(\mem<13><15> ), .B(n1251), .Y(n1615) );
  OAI21X1 U1448 ( .A(n126), .B(n1293), .C(n1615), .Y(n2041) );
  NAND2X1 U1449 ( .A(\mem<12><0> ), .B(n1252), .Y(n1616) );
  OAI21X1 U1450 ( .A(n128), .B(n1270), .C(n1616), .Y(n2040) );
  NAND2X1 U1451 ( .A(\mem<12><1> ), .B(n1252), .Y(n1617) );
  OAI21X1 U1452 ( .A(n128), .B(n1272), .C(n1617), .Y(n2039) );
  NAND2X1 U1453 ( .A(\mem<12><2> ), .B(n1252), .Y(n1618) );
  OAI21X1 U1454 ( .A(n128), .B(n1273), .C(n1618), .Y(n2038) );
  NAND2X1 U1455 ( .A(\mem<12><3> ), .B(n1252), .Y(n1619) );
  OAI21X1 U1456 ( .A(n128), .B(n1274), .C(n1619), .Y(n2037) );
  NAND2X1 U1457 ( .A(\mem<12><4> ), .B(n1252), .Y(n1620) );
  OAI21X1 U1458 ( .A(n128), .B(n1275), .C(n1620), .Y(n2036) );
  NAND2X1 U1459 ( .A(\mem<12><5> ), .B(n1252), .Y(n1621) );
  OAI21X1 U1460 ( .A(n128), .B(n1277), .C(n1621), .Y(n2035) );
  NAND2X1 U1461 ( .A(\mem<12><6> ), .B(n1252), .Y(n1622) );
  OAI21X1 U1462 ( .A(n128), .B(n1278), .C(n1622), .Y(n2034) );
  NAND2X1 U1463 ( .A(\mem<12><7> ), .B(n1252), .Y(n1623) );
  OAI21X1 U1464 ( .A(n128), .B(n1279), .C(n1623), .Y(n2033) );
  NAND2X1 U1465 ( .A(\mem<12><8> ), .B(n1253), .Y(n1624) );
  OAI21X1 U1466 ( .A(n128), .B(n1280), .C(n1624), .Y(n2032) );
  NAND2X1 U1467 ( .A(\mem<12><9> ), .B(n1253), .Y(n1625) );
  OAI21X1 U1468 ( .A(n128), .B(n1282), .C(n1625), .Y(n2031) );
  NAND2X1 U1469 ( .A(\mem<12><10> ), .B(n1253), .Y(n1626) );
  OAI21X1 U1470 ( .A(n128), .B(n1283), .C(n1626), .Y(n2030) );
  NAND2X1 U1471 ( .A(\mem<12><11> ), .B(n1253), .Y(n1627) );
  OAI21X1 U1472 ( .A(n128), .B(n1285), .C(n1627), .Y(n2029) );
  NAND2X1 U1473 ( .A(\mem<12><12> ), .B(n1253), .Y(n1628) );
  OAI21X1 U1474 ( .A(n128), .B(n1287), .C(n1628), .Y(n2028) );
  NAND2X1 U1475 ( .A(\mem<12><13> ), .B(n1253), .Y(n1629) );
  OAI21X1 U1476 ( .A(n128), .B(n1289), .C(n1629), .Y(n2027) );
  NAND2X1 U1477 ( .A(\mem<12><14> ), .B(n1253), .Y(n1630) );
  OAI21X1 U1478 ( .A(n128), .B(n1291), .C(n1630), .Y(n2026) );
  NAND2X1 U1479 ( .A(\mem<12><15> ), .B(n1253), .Y(n1631) );
  OAI21X1 U1480 ( .A(n128), .B(n1293), .C(n1631), .Y(n2025) );
  NAND2X1 U1481 ( .A(\mem<11><0> ), .B(n1254), .Y(n1632) );
  OAI21X1 U1482 ( .A(n130), .B(n1270), .C(n1632), .Y(n2024) );
  NAND2X1 U1483 ( .A(\mem<11><1> ), .B(n1254), .Y(n1633) );
  OAI21X1 U1484 ( .A(n130), .B(n1271), .C(n1633), .Y(n2023) );
  NAND2X1 U1485 ( .A(\mem<11><2> ), .B(n1254), .Y(n1634) );
  OAI21X1 U1486 ( .A(n130), .B(n1273), .C(n1634), .Y(n2022) );
  NAND2X1 U1487 ( .A(\mem<11><3> ), .B(n1254), .Y(n1635) );
  OAI21X1 U1488 ( .A(n130), .B(n1274), .C(n1635), .Y(n2021) );
  NAND2X1 U1489 ( .A(\mem<11><4> ), .B(n1254), .Y(n1636) );
  OAI21X1 U1490 ( .A(n130), .B(n1275), .C(n1636), .Y(n2020) );
  NAND2X1 U1491 ( .A(\mem<11><5> ), .B(n1254), .Y(n1637) );
  OAI21X1 U1492 ( .A(n130), .B(n1276), .C(n1637), .Y(n2019) );
  NAND2X1 U1493 ( .A(\mem<11><6> ), .B(n1254), .Y(n1638) );
  OAI21X1 U1494 ( .A(n130), .B(n1278), .C(n1638), .Y(n2018) );
  NAND2X1 U1495 ( .A(\mem<11><7> ), .B(n1254), .Y(n1639) );
  OAI21X1 U1496 ( .A(n130), .B(n1279), .C(n1639), .Y(n2017) );
  NAND2X1 U1497 ( .A(\mem<11><8> ), .B(n1255), .Y(n1640) );
  OAI21X1 U1498 ( .A(n130), .B(n1280), .C(n1640), .Y(n2016) );
  NAND2X1 U1499 ( .A(\mem<11><9> ), .B(n1255), .Y(n1641) );
  OAI21X1 U1500 ( .A(n130), .B(n1281), .C(n1641), .Y(n2015) );
  NAND2X1 U1501 ( .A(\mem<11><10> ), .B(n1255), .Y(n1642) );
  OAI21X1 U1502 ( .A(n130), .B(n1283), .C(n1642), .Y(n2014) );
  NAND2X1 U1503 ( .A(\mem<11><11> ), .B(n1255), .Y(n1643) );
  OAI21X1 U1504 ( .A(n130), .B(n1284), .C(n1643), .Y(n2013) );
  NAND2X1 U1505 ( .A(\mem<11><12> ), .B(n1255), .Y(n1644) );
  OAI21X1 U1506 ( .A(n130), .B(n1286), .C(n1644), .Y(n2012) );
  NAND2X1 U1507 ( .A(\mem<11><13> ), .B(n1255), .Y(n1645) );
  OAI21X1 U1508 ( .A(n130), .B(n1288), .C(n1645), .Y(n2011) );
  NAND2X1 U1509 ( .A(\mem<11><14> ), .B(n1255), .Y(n1646) );
  OAI21X1 U1510 ( .A(n130), .B(n1290), .C(n1646), .Y(n2010) );
  NAND2X1 U1511 ( .A(\mem<11><15> ), .B(n1255), .Y(n1647) );
  OAI21X1 U1512 ( .A(n130), .B(n1292), .C(n1647), .Y(n2009) );
  NAND2X1 U1513 ( .A(\mem<10><0> ), .B(n1256), .Y(n1648) );
  OAI21X1 U1514 ( .A(n132), .B(n1270), .C(n1648), .Y(n2008) );
  NAND2X1 U1515 ( .A(\mem<10><1> ), .B(n1256), .Y(n1649) );
  OAI21X1 U1516 ( .A(n132), .B(n1271), .C(n1649), .Y(n2007) );
  NAND2X1 U1517 ( .A(\mem<10><2> ), .B(n1256), .Y(n1650) );
  OAI21X1 U1518 ( .A(n132), .B(n1273), .C(n1650), .Y(n2006) );
  NAND2X1 U1519 ( .A(\mem<10><3> ), .B(n1256), .Y(n1651) );
  OAI21X1 U1520 ( .A(n132), .B(n1274), .C(n1651), .Y(n2005) );
  NAND2X1 U1521 ( .A(\mem<10><4> ), .B(n1256), .Y(n1652) );
  OAI21X1 U1522 ( .A(n132), .B(n1275), .C(n1652), .Y(n2004) );
  NAND2X1 U1523 ( .A(\mem<10><5> ), .B(n1256), .Y(n1653) );
  OAI21X1 U1524 ( .A(n132), .B(n1276), .C(n1653), .Y(n2003) );
  NAND2X1 U1525 ( .A(\mem<10><6> ), .B(n1256), .Y(n1654) );
  OAI21X1 U1526 ( .A(n132), .B(n1278), .C(n1654), .Y(n2002) );
  NAND2X1 U1527 ( .A(\mem<10><7> ), .B(n1256), .Y(n1655) );
  OAI21X1 U1528 ( .A(n132), .B(n1279), .C(n1655), .Y(n2001) );
  NAND2X1 U1529 ( .A(\mem<10><8> ), .B(n1257), .Y(n1656) );
  OAI21X1 U1530 ( .A(n132), .B(n1280), .C(n1656), .Y(n2000) );
  NAND2X1 U1531 ( .A(\mem<10><9> ), .B(n1257), .Y(n1657) );
  OAI21X1 U1532 ( .A(n132), .B(n1281), .C(n1657), .Y(n1999) );
  NAND2X1 U1533 ( .A(\mem<10><10> ), .B(n1257), .Y(n1658) );
  OAI21X1 U1534 ( .A(n132), .B(n1283), .C(n1658), .Y(n1998) );
  NAND2X1 U1535 ( .A(\mem<10><11> ), .B(n1257), .Y(n1659) );
  OAI21X1 U1536 ( .A(n132), .B(n1284), .C(n1659), .Y(n1997) );
  NAND2X1 U1537 ( .A(\mem<10><12> ), .B(n1257), .Y(n1660) );
  OAI21X1 U1538 ( .A(n132), .B(n1286), .C(n1660), .Y(n1996) );
  NAND2X1 U1539 ( .A(\mem<10><13> ), .B(n1257), .Y(n1661) );
  OAI21X1 U1540 ( .A(n132), .B(n1288), .C(n1661), .Y(n1995) );
  NAND2X1 U1541 ( .A(\mem<10><14> ), .B(n1257), .Y(n1662) );
  OAI21X1 U1542 ( .A(n132), .B(n1290), .C(n1662), .Y(n1994) );
  NAND2X1 U1543 ( .A(\mem<10><15> ), .B(n1257), .Y(n1663) );
  OAI21X1 U1544 ( .A(n132), .B(n1292), .C(n1663), .Y(n1993) );
  NAND2X1 U1545 ( .A(\mem<9><0> ), .B(n1258), .Y(n1664) );
  OAI21X1 U1546 ( .A(n134), .B(n1270), .C(n1664), .Y(n1992) );
  NAND2X1 U1547 ( .A(\mem<9><1> ), .B(n1258), .Y(n1665) );
  OAI21X1 U1548 ( .A(n134), .B(n1271), .C(n1665), .Y(n1991) );
  NAND2X1 U1549 ( .A(\mem<9><2> ), .B(n1258), .Y(n1666) );
  OAI21X1 U1550 ( .A(n134), .B(n1273), .C(n1666), .Y(n1990) );
  NAND2X1 U1551 ( .A(\mem<9><3> ), .B(n1258), .Y(n1667) );
  OAI21X1 U1552 ( .A(n134), .B(n1274), .C(n1667), .Y(n1989) );
  NAND2X1 U1553 ( .A(\mem<9><4> ), .B(n1258), .Y(n1668) );
  OAI21X1 U1554 ( .A(n134), .B(n1275), .C(n1668), .Y(n1988) );
  NAND2X1 U1555 ( .A(\mem<9><5> ), .B(n1258), .Y(n1669) );
  OAI21X1 U1556 ( .A(n134), .B(n1276), .C(n1669), .Y(n1987) );
  NAND2X1 U1557 ( .A(\mem<9><6> ), .B(n1258), .Y(n1670) );
  OAI21X1 U1558 ( .A(n134), .B(n1278), .C(n1670), .Y(n1986) );
  NAND2X1 U1559 ( .A(\mem<9><7> ), .B(n1258), .Y(n1671) );
  OAI21X1 U1560 ( .A(n134), .B(n1279), .C(n1671), .Y(n1985) );
  NAND2X1 U1561 ( .A(\mem<9><8> ), .B(n1259), .Y(n1672) );
  OAI21X1 U1562 ( .A(n134), .B(n1280), .C(n1672), .Y(n1984) );
  NAND2X1 U1563 ( .A(\mem<9><9> ), .B(n1259), .Y(n1673) );
  OAI21X1 U1564 ( .A(n134), .B(n1281), .C(n1673), .Y(n1983) );
  NAND2X1 U1565 ( .A(\mem<9><10> ), .B(n1259), .Y(n1674) );
  OAI21X1 U1566 ( .A(n134), .B(n1283), .C(n1674), .Y(n1982) );
  NAND2X1 U1567 ( .A(\mem<9><11> ), .B(n1259), .Y(n1675) );
  OAI21X1 U1568 ( .A(n134), .B(n1284), .C(n1675), .Y(n1981) );
  NAND2X1 U1569 ( .A(\mem<9><12> ), .B(n1259), .Y(n1676) );
  OAI21X1 U1570 ( .A(n134), .B(n1286), .C(n1676), .Y(n1980) );
  NAND2X1 U1571 ( .A(\mem<9><13> ), .B(n1259), .Y(n1677) );
  OAI21X1 U1572 ( .A(n134), .B(n1288), .C(n1677), .Y(n1979) );
  NAND2X1 U1573 ( .A(\mem<9><14> ), .B(n1259), .Y(n1678) );
  OAI21X1 U1574 ( .A(n134), .B(n1290), .C(n1678), .Y(n1978) );
  NAND2X1 U1575 ( .A(\mem<9><15> ), .B(n1259), .Y(n1679) );
  OAI21X1 U1576 ( .A(n134), .B(n1292), .C(n1679), .Y(n1977) );
  NAND2X1 U1577 ( .A(\mem<8><0> ), .B(n1261), .Y(n1681) );
  OAI21X1 U1578 ( .A(n1260), .B(n1270), .C(n1681), .Y(n1976) );
  NAND2X1 U1579 ( .A(\mem<8><1> ), .B(n1261), .Y(n1682) );
  OAI21X1 U1580 ( .A(n1260), .B(n1271), .C(n1682), .Y(n1975) );
  NAND2X1 U1581 ( .A(\mem<8><2> ), .B(n1261), .Y(n1683) );
  OAI21X1 U1582 ( .A(n1260), .B(n1273), .C(n1683), .Y(n1974) );
  NAND2X1 U1583 ( .A(\mem<8><3> ), .B(n1261), .Y(n1684) );
  OAI21X1 U1584 ( .A(n1260), .B(n1274), .C(n1684), .Y(n1973) );
  NAND2X1 U1585 ( .A(\mem<8><4> ), .B(n1261), .Y(n1685) );
  OAI21X1 U1586 ( .A(n1260), .B(n1275), .C(n1685), .Y(n1972) );
  NAND2X1 U1587 ( .A(\mem<8><5> ), .B(n1261), .Y(n1686) );
  OAI21X1 U1588 ( .A(n1260), .B(n1276), .C(n1686), .Y(n1971) );
  NAND2X1 U1589 ( .A(\mem<8><6> ), .B(n1261), .Y(n1687) );
  OAI21X1 U1590 ( .A(n1260), .B(n1278), .C(n1687), .Y(n1970) );
  NAND2X1 U1591 ( .A(\mem<8><7> ), .B(n1261), .Y(n1688) );
  OAI21X1 U1592 ( .A(n1260), .B(n1279), .C(n1688), .Y(n1969) );
  NAND2X1 U1593 ( .A(\mem<8><8> ), .B(n1262), .Y(n1689) );
  OAI21X1 U1594 ( .A(n1260), .B(n1280), .C(n1689), .Y(n1968) );
  NAND2X1 U1595 ( .A(\mem<8><9> ), .B(n1262), .Y(n1690) );
  OAI21X1 U1596 ( .A(n1260), .B(n1281), .C(n1690), .Y(n1967) );
  NAND2X1 U1597 ( .A(\mem<8><10> ), .B(n1262), .Y(n1691) );
  OAI21X1 U1598 ( .A(n1260), .B(n1283), .C(n1691), .Y(n1966) );
  NAND2X1 U1599 ( .A(\mem<8><11> ), .B(n1262), .Y(n1692) );
  OAI21X1 U1600 ( .A(n1260), .B(n1284), .C(n1692), .Y(n1965) );
  NAND2X1 U1601 ( .A(\mem<8><12> ), .B(n1262), .Y(n1693) );
  OAI21X1 U1602 ( .A(n1260), .B(n1286), .C(n1693), .Y(n1964) );
  NAND2X1 U1603 ( .A(\mem<8><13> ), .B(n1262), .Y(n1694) );
  OAI21X1 U1604 ( .A(n1260), .B(n1288), .C(n1694), .Y(n1963) );
  NAND2X1 U1605 ( .A(\mem<8><14> ), .B(n1262), .Y(n1695) );
  OAI21X1 U1606 ( .A(n1260), .B(n1290), .C(n1695), .Y(n1962) );
  NAND2X1 U1607 ( .A(\mem<8><15> ), .B(n1262), .Y(n1696) );
  OAI21X1 U1608 ( .A(n1260), .B(n1292), .C(n1696), .Y(n1961) );
  NAND3X1 U1609 ( .A(n1301), .B(n2345), .C(n1303), .Y(n1697) );
  NAND2X1 U1610 ( .A(\mem<7><0> ), .B(n137), .Y(n1698) );
  OAI21X1 U1611 ( .A(n136), .B(n1270), .C(n1698), .Y(n1960) );
  NAND2X1 U1612 ( .A(\mem<7><1> ), .B(n137), .Y(n1699) );
  OAI21X1 U1613 ( .A(n136), .B(n1271), .C(n1699), .Y(n1959) );
  NAND2X1 U1614 ( .A(\mem<7><2> ), .B(n137), .Y(n1700) );
  OAI21X1 U1615 ( .A(n136), .B(n1273), .C(n1700), .Y(n1958) );
  NAND2X1 U1616 ( .A(\mem<7><3> ), .B(n137), .Y(n1701) );
  OAI21X1 U1617 ( .A(n136), .B(n1274), .C(n1701), .Y(n1957) );
  NAND2X1 U1618 ( .A(\mem<7><4> ), .B(n137), .Y(n1702) );
  OAI21X1 U1619 ( .A(n136), .B(n1275), .C(n1702), .Y(n1956) );
  NAND2X1 U1620 ( .A(\mem<7><5> ), .B(n137), .Y(n1703) );
  OAI21X1 U1621 ( .A(n136), .B(n1276), .C(n1703), .Y(n1955) );
  NAND2X1 U1622 ( .A(\mem<7><6> ), .B(n137), .Y(n1704) );
  OAI21X1 U1623 ( .A(n136), .B(n1278), .C(n1704), .Y(n1954) );
  NAND2X1 U1624 ( .A(\mem<7><7> ), .B(n137), .Y(n1705) );
  OAI21X1 U1625 ( .A(n136), .B(n1279), .C(n1705), .Y(n1953) );
  NAND2X1 U1626 ( .A(\mem<7><8> ), .B(n137), .Y(n1706) );
  OAI21X1 U1627 ( .A(n136), .B(n1280), .C(n1706), .Y(n1952) );
  NAND2X1 U1628 ( .A(\mem<7><9> ), .B(n137), .Y(n1707) );
  OAI21X1 U1629 ( .A(n136), .B(n1281), .C(n1707), .Y(n1951) );
  NAND2X1 U1630 ( .A(\mem<7><10> ), .B(n137), .Y(n1708) );
  OAI21X1 U1631 ( .A(n136), .B(n1283), .C(n1708), .Y(n1950) );
  NAND2X1 U1632 ( .A(\mem<7><11> ), .B(n137), .Y(n1709) );
  OAI21X1 U1633 ( .A(n136), .B(n1284), .C(n1709), .Y(n1949) );
  NAND2X1 U1634 ( .A(\mem<7><12> ), .B(n137), .Y(n1710) );
  OAI21X1 U1635 ( .A(n136), .B(n1286), .C(n1710), .Y(n1948) );
  NAND2X1 U1636 ( .A(\mem<7><13> ), .B(n137), .Y(n1711) );
  OAI21X1 U1637 ( .A(n136), .B(n1288), .C(n1711), .Y(n1947) );
  NAND2X1 U1638 ( .A(\mem<7><14> ), .B(n137), .Y(n1712) );
  OAI21X1 U1639 ( .A(n136), .B(n1290), .C(n1712), .Y(n1946) );
  NAND2X1 U1640 ( .A(\mem<7><15> ), .B(n137), .Y(n1713) );
  OAI21X1 U1641 ( .A(n136), .B(n1292), .C(n1713), .Y(n1945) );
  NAND2X1 U1642 ( .A(\mem<6><0> ), .B(n140), .Y(n1714) );
  OAI21X1 U1643 ( .A(n139), .B(n1270), .C(n1714), .Y(n1944) );
  NAND2X1 U1644 ( .A(\mem<6><1> ), .B(n140), .Y(n1715) );
  OAI21X1 U1645 ( .A(n139), .B(n1271), .C(n1715), .Y(n1943) );
  NAND2X1 U1646 ( .A(\mem<6><2> ), .B(n140), .Y(n1716) );
  OAI21X1 U1647 ( .A(n139), .B(n1273), .C(n1716), .Y(n1942) );
  NAND2X1 U1648 ( .A(\mem<6><3> ), .B(n140), .Y(n1717) );
  OAI21X1 U1649 ( .A(n139), .B(n1274), .C(n1717), .Y(n1941) );
  NAND2X1 U1650 ( .A(\mem<6><4> ), .B(n140), .Y(n1718) );
  OAI21X1 U1651 ( .A(n139), .B(n1275), .C(n1718), .Y(n1940) );
  NAND2X1 U1652 ( .A(\mem<6><5> ), .B(n140), .Y(n1719) );
  OAI21X1 U1653 ( .A(n139), .B(n1276), .C(n1719), .Y(n1939) );
  NAND2X1 U1654 ( .A(\mem<6><6> ), .B(n140), .Y(n1720) );
  OAI21X1 U1655 ( .A(n139), .B(n1278), .C(n1720), .Y(n1938) );
  NAND2X1 U1656 ( .A(\mem<6><7> ), .B(n140), .Y(n1721) );
  OAI21X1 U1657 ( .A(n139), .B(n1279), .C(n1721), .Y(n1937) );
  NAND2X1 U1658 ( .A(\mem<6><8> ), .B(n140), .Y(n1722) );
  OAI21X1 U1659 ( .A(n139), .B(n1280), .C(n1722), .Y(n1936) );
  NAND2X1 U1660 ( .A(\mem<6><9> ), .B(n140), .Y(n1723) );
  OAI21X1 U1661 ( .A(n139), .B(n1281), .C(n1723), .Y(n1935) );
  NAND2X1 U1662 ( .A(\mem<6><10> ), .B(n140), .Y(n1724) );
  OAI21X1 U1663 ( .A(n139), .B(n1283), .C(n1724), .Y(n1934) );
  NAND2X1 U1664 ( .A(\mem<6><11> ), .B(n140), .Y(n1725) );
  OAI21X1 U1665 ( .A(n139), .B(n1284), .C(n1725), .Y(n1933) );
  NAND2X1 U1666 ( .A(\mem<6><12> ), .B(n140), .Y(n1726) );
  OAI21X1 U1667 ( .A(n139), .B(n1286), .C(n1726), .Y(n1932) );
  NAND2X1 U1668 ( .A(\mem<6><13> ), .B(n140), .Y(n1727) );
  OAI21X1 U1669 ( .A(n139), .B(n1288), .C(n1727), .Y(n1931) );
  NAND2X1 U1670 ( .A(\mem<6><14> ), .B(n140), .Y(n1728) );
  OAI21X1 U1671 ( .A(n139), .B(n1290), .C(n1728), .Y(n1930) );
  NAND2X1 U1672 ( .A(\mem<6><15> ), .B(n140), .Y(n1729) );
  OAI21X1 U1673 ( .A(n139), .B(n1292), .C(n1729), .Y(n1929) );
  NAND2X1 U1674 ( .A(\mem<5><0> ), .B(n144), .Y(n1731) );
  OAI21X1 U1675 ( .A(n142), .B(n1270), .C(n1731), .Y(n1928) );
  NAND2X1 U1676 ( .A(\mem<5><1> ), .B(n144), .Y(n1732) );
  OAI21X1 U1677 ( .A(n142), .B(n1271), .C(n1732), .Y(n1927) );
  NAND2X1 U1678 ( .A(\mem<5><2> ), .B(n144), .Y(n1733) );
  OAI21X1 U1679 ( .A(n142), .B(n1273), .C(n1733), .Y(n1926) );
  NAND2X1 U1680 ( .A(\mem<5><3> ), .B(n144), .Y(n1734) );
  OAI21X1 U1681 ( .A(n142), .B(n1274), .C(n1734), .Y(n1925) );
  NAND2X1 U1682 ( .A(\mem<5><4> ), .B(n144), .Y(n1735) );
  OAI21X1 U1683 ( .A(n142), .B(n1275), .C(n1735), .Y(n1924) );
  NAND2X1 U1684 ( .A(\mem<5><5> ), .B(n144), .Y(n1736) );
  OAI21X1 U1685 ( .A(n142), .B(n1276), .C(n1736), .Y(n1923) );
  NAND2X1 U1686 ( .A(\mem<5><6> ), .B(n144), .Y(n1737) );
  OAI21X1 U1687 ( .A(n142), .B(n1278), .C(n1737), .Y(n1922) );
  NAND2X1 U1688 ( .A(\mem<5><7> ), .B(n144), .Y(n1738) );
  OAI21X1 U1689 ( .A(n142), .B(n1279), .C(n1738), .Y(n1921) );
  NAND2X1 U1690 ( .A(\mem<5><8> ), .B(n143), .Y(n1739) );
  OAI21X1 U1691 ( .A(n142), .B(n1280), .C(n1739), .Y(n1920) );
  NAND2X1 U1692 ( .A(\mem<5><9> ), .B(n143), .Y(n1740) );
  OAI21X1 U1693 ( .A(n142), .B(n1281), .C(n1740), .Y(n1919) );
  NAND2X1 U1694 ( .A(\mem<5><10> ), .B(n143), .Y(n1741) );
  OAI21X1 U1695 ( .A(n142), .B(n1283), .C(n1741), .Y(n1918) );
  NAND2X1 U1696 ( .A(\mem<5><11> ), .B(n143), .Y(n1742) );
  OAI21X1 U1697 ( .A(n142), .B(n1284), .C(n1742), .Y(n1917) );
  NAND2X1 U1698 ( .A(\mem<5><12> ), .B(n143), .Y(n1743) );
  OAI21X1 U1699 ( .A(n142), .B(n1286), .C(n1743), .Y(n1916) );
  NAND2X1 U1700 ( .A(\mem<5><13> ), .B(n143), .Y(n1744) );
  OAI21X1 U1701 ( .A(n142), .B(n1288), .C(n1744), .Y(n1915) );
  NAND2X1 U1702 ( .A(\mem<5><14> ), .B(n143), .Y(n1745) );
  OAI21X1 U1703 ( .A(n142), .B(n1290), .C(n1745), .Y(n1914) );
  NAND2X1 U1704 ( .A(\mem<5><15> ), .B(n143), .Y(n1746) );
  OAI21X1 U1705 ( .A(n142), .B(n1292), .C(n1746), .Y(n1913) );
  NAND2X1 U1706 ( .A(\mem<4><0> ), .B(n148), .Y(n1748) );
  OAI21X1 U1707 ( .A(n146), .B(n1270), .C(n1748), .Y(n1912) );
  NAND2X1 U1708 ( .A(\mem<4><1> ), .B(n148), .Y(n1749) );
  OAI21X1 U1709 ( .A(n146), .B(n1271), .C(n1749), .Y(n1911) );
  NAND2X1 U1710 ( .A(\mem<4><2> ), .B(n148), .Y(n1750) );
  OAI21X1 U1711 ( .A(n146), .B(n1273), .C(n1750), .Y(n1910) );
  NAND2X1 U1712 ( .A(\mem<4><3> ), .B(n148), .Y(n1751) );
  OAI21X1 U1713 ( .A(n146), .B(n1274), .C(n1751), .Y(n1909) );
  NAND2X1 U1714 ( .A(\mem<4><4> ), .B(n148), .Y(n1752) );
  OAI21X1 U1715 ( .A(n146), .B(n1275), .C(n1752), .Y(n1908) );
  NAND2X1 U1716 ( .A(\mem<4><5> ), .B(n148), .Y(n1753) );
  OAI21X1 U1717 ( .A(n146), .B(n1276), .C(n1753), .Y(n1907) );
  NAND2X1 U1718 ( .A(\mem<4><6> ), .B(n148), .Y(n1754) );
  OAI21X1 U1719 ( .A(n146), .B(n1278), .C(n1754), .Y(n1906) );
  NAND2X1 U1720 ( .A(\mem<4><7> ), .B(n148), .Y(n1755) );
  OAI21X1 U1721 ( .A(n146), .B(n1279), .C(n1755), .Y(n1905) );
  NAND2X1 U1722 ( .A(\mem<4><8> ), .B(n147), .Y(n1756) );
  OAI21X1 U1723 ( .A(n146), .B(n1280), .C(n1756), .Y(n1904) );
  NAND2X1 U1724 ( .A(\mem<4><9> ), .B(n147), .Y(n1757) );
  OAI21X1 U1725 ( .A(n146), .B(n1281), .C(n1757), .Y(n1903) );
  NAND2X1 U1726 ( .A(\mem<4><10> ), .B(n147), .Y(n1758) );
  OAI21X1 U1727 ( .A(n146), .B(n1283), .C(n1758), .Y(n1902) );
  NAND2X1 U1728 ( .A(\mem<4><11> ), .B(n147), .Y(n1759) );
  OAI21X1 U1729 ( .A(n146), .B(n1284), .C(n1759), .Y(n1901) );
  NAND2X1 U1730 ( .A(\mem<4><12> ), .B(n147), .Y(n1760) );
  OAI21X1 U1731 ( .A(n146), .B(n1286), .C(n1760), .Y(n1900) );
  NAND2X1 U1732 ( .A(\mem<4><13> ), .B(n147), .Y(n1761) );
  OAI21X1 U1733 ( .A(n146), .B(n1288), .C(n1761), .Y(n1899) );
  NAND2X1 U1734 ( .A(\mem<4><14> ), .B(n147), .Y(n1762) );
  OAI21X1 U1735 ( .A(n146), .B(n1290), .C(n1762), .Y(n1898) );
  NAND2X1 U1736 ( .A(\mem<4><15> ), .B(n147), .Y(n1763) );
  OAI21X1 U1737 ( .A(n146), .B(n1292), .C(n1763), .Y(n1897) );
  NAND2X1 U1738 ( .A(\mem<3><0> ), .B(n152), .Y(n1765) );
  OAI21X1 U1739 ( .A(n150), .B(n1270), .C(n1765), .Y(n1896) );
  NAND2X1 U1740 ( .A(\mem<3><1> ), .B(n152), .Y(n1766) );
  OAI21X1 U1741 ( .A(n150), .B(n1271), .C(n1766), .Y(n1895) );
  NAND2X1 U1742 ( .A(\mem<3><2> ), .B(n152), .Y(n1767) );
  OAI21X1 U1743 ( .A(n150), .B(n1273), .C(n1767), .Y(n1894) );
  NAND2X1 U1744 ( .A(\mem<3><3> ), .B(n152), .Y(n1768) );
  OAI21X1 U1745 ( .A(n150), .B(n1274), .C(n1768), .Y(n1893) );
  NAND2X1 U1746 ( .A(\mem<3><4> ), .B(n152), .Y(n1769) );
  OAI21X1 U1747 ( .A(n150), .B(n1275), .C(n1769), .Y(n1892) );
  NAND2X1 U1748 ( .A(\mem<3><5> ), .B(n152), .Y(n1770) );
  OAI21X1 U1749 ( .A(n150), .B(n1276), .C(n1770), .Y(n1891) );
  NAND2X1 U1750 ( .A(\mem<3><6> ), .B(n152), .Y(n1771) );
  OAI21X1 U1751 ( .A(n150), .B(n1278), .C(n1771), .Y(n1890) );
  NAND2X1 U1752 ( .A(\mem<3><7> ), .B(n152), .Y(n1772) );
  OAI21X1 U1753 ( .A(n150), .B(n1279), .C(n1772), .Y(n1889) );
  NAND2X1 U1754 ( .A(\mem<3><8> ), .B(n151), .Y(n1773) );
  OAI21X1 U1755 ( .A(n150), .B(n1280), .C(n1773), .Y(n1888) );
  NAND2X1 U1756 ( .A(\mem<3><9> ), .B(n151), .Y(n1774) );
  OAI21X1 U1757 ( .A(n150), .B(n1281), .C(n1774), .Y(n1887) );
  NAND2X1 U1758 ( .A(\mem<3><10> ), .B(n151), .Y(n1775) );
  OAI21X1 U1759 ( .A(n150), .B(n1283), .C(n1775), .Y(n1886) );
  NAND2X1 U1760 ( .A(\mem<3><11> ), .B(n151), .Y(n1776) );
  OAI21X1 U1761 ( .A(n150), .B(n1284), .C(n1776), .Y(n1885) );
  NAND2X1 U1762 ( .A(\mem<3><12> ), .B(n151), .Y(n1777) );
  OAI21X1 U1763 ( .A(n150), .B(n1286), .C(n1777), .Y(n1884) );
  NAND2X1 U1764 ( .A(\mem<3><13> ), .B(n151), .Y(n1778) );
  OAI21X1 U1765 ( .A(n150), .B(n1288), .C(n1778), .Y(n1883) );
  NAND2X1 U1766 ( .A(\mem<3><14> ), .B(n151), .Y(n1779) );
  OAI21X1 U1767 ( .A(n150), .B(n1290), .C(n1779), .Y(n1882) );
  NAND2X1 U1768 ( .A(\mem<3><15> ), .B(n151), .Y(n1780) );
  OAI21X1 U1769 ( .A(n150), .B(n1292), .C(n1780), .Y(n1881) );
  NAND2X1 U1770 ( .A(\mem<2><0> ), .B(n156), .Y(n1782) );
  OAI21X1 U1771 ( .A(n154), .B(n1270), .C(n1782), .Y(n1880) );
  NAND2X1 U1772 ( .A(\mem<2><1> ), .B(n156), .Y(n1783) );
  OAI21X1 U1773 ( .A(n154), .B(n1271), .C(n1783), .Y(n1879) );
  NAND2X1 U1774 ( .A(\mem<2><2> ), .B(n156), .Y(n1784) );
  OAI21X1 U1775 ( .A(n154), .B(n1273), .C(n1784), .Y(n1878) );
  NAND2X1 U1776 ( .A(\mem<2><3> ), .B(n156), .Y(n1785) );
  OAI21X1 U1777 ( .A(n154), .B(n1274), .C(n1785), .Y(n1877) );
  NAND2X1 U1778 ( .A(\mem<2><4> ), .B(n156), .Y(n1786) );
  OAI21X1 U1779 ( .A(n154), .B(n1275), .C(n1786), .Y(n1876) );
  NAND2X1 U1780 ( .A(\mem<2><5> ), .B(n156), .Y(n1787) );
  OAI21X1 U1781 ( .A(n154), .B(n1276), .C(n1787), .Y(n1875) );
  NAND2X1 U1782 ( .A(\mem<2><6> ), .B(n156), .Y(n1788) );
  OAI21X1 U1783 ( .A(n154), .B(n1278), .C(n1788), .Y(n1874) );
  NAND2X1 U1784 ( .A(\mem<2><7> ), .B(n156), .Y(n1789) );
  OAI21X1 U1785 ( .A(n154), .B(n1279), .C(n1789), .Y(n1873) );
  NAND2X1 U1786 ( .A(\mem<2><8> ), .B(n155), .Y(n1790) );
  OAI21X1 U1787 ( .A(n154), .B(n1280), .C(n1790), .Y(n1872) );
  NAND2X1 U1788 ( .A(\mem<2><9> ), .B(n155), .Y(n1791) );
  OAI21X1 U1789 ( .A(n154), .B(n1281), .C(n1791), .Y(n1871) );
  NAND2X1 U1790 ( .A(\mem<2><10> ), .B(n155), .Y(n1792) );
  OAI21X1 U1791 ( .A(n154), .B(n1283), .C(n1792), .Y(n1870) );
  NAND2X1 U1792 ( .A(\mem<2><11> ), .B(n155), .Y(n1793) );
  OAI21X1 U1793 ( .A(n154), .B(n1284), .C(n1793), .Y(n1869) );
  NAND2X1 U1794 ( .A(\mem<2><12> ), .B(n155), .Y(n1794) );
  OAI21X1 U1795 ( .A(n154), .B(n1286), .C(n1794), .Y(n1868) );
  NAND2X1 U1796 ( .A(\mem<2><13> ), .B(n155), .Y(n1795) );
  OAI21X1 U1797 ( .A(n154), .B(n1288), .C(n1795), .Y(n1867) );
  NAND2X1 U1798 ( .A(\mem<2><14> ), .B(n155), .Y(n1796) );
  OAI21X1 U1799 ( .A(n154), .B(n1290), .C(n1796), .Y(n1866) );
  NAND2X1 U1800 ( .A(\mem<2><15> ), .B(n155), .Y(n1797) );
  OAI21X1 U1801 ( .A(n154), .B(n1292), .C(n1797), .Y(n1865) );
  NAND2X1 U1802 ( .A(\mem<1><0> ), .B(n160), .Y(n1799) );
  OAI21X1 U1803 ( .A(n158), .B(n1270), .C(n1799), .Y(n1864) );
  NAND2X1 U1804 ( .A(\mem<1><1> ), .B(n160), .Y(n1800) );
  OAI21X1 U1805 ( .A(n158), .B(n1271), .C(n1800), .Y(n1863) );
  NAND2X1 U1806 ( .A(\mem<1><2> ), .B(n160), .Y(n1801) );
  OAI21X1 U1807 ( .A(n158), .B(n1273), .C(n1801), .Y(n1862) );
  NAND2X1 U1808 ( .A(\mem<1><3> ), .B(n160), .Y(n1802) );
  OAI21X1 U1809 ( .A(n158), .B(n1274), .C(n1802), .Y(n1861) );
  NAND2X1 U1810 ( .A(\mem<1><4> ), .B(n160), .Y(n1803) );
  OAI21X1 U1811 ( .A(n158), .B(n1275), .C(n1803), .Y(n1860) );
  NAND2X1 U1812 ( .A(\mem<1><5> ), .B(n160), .Y(n1804) );
  OAI21X1 U1813 ( .A(n158), .B(n1276), .C(n1804), .Y(n1859) );
  NAND2X1 U1814 ( .A(\mem<1><6> ), .B(n160), .Y(n1805) );
  OAI21X1 U1815 ( .A(n158), .B(n1278), .C(n1805), .Y(n1858) );
  NAND2X1 U1816 ( .A(\mem<1><7> ), .B(n160), .Y(n1806) );
  OAI21X1 U1817 ( .A(n158), .B(n1279), .C(n1806), .Y(n1857) );
  NAND2X1 U1818 ( .A(\mem<1><8> ), .B(n159), .Y(n1807) );
  OAI21X1 U1819 ( .A(n158), .B(n1280), .C(n1807), .Y(n1856) );
  NAND2X1 U1820 ( .A(\mem<1><9> ), .B(n159), .Y(n1808) );
  OAI21X1 U1821 ( .A(n158), .B(n1281), .C(n1808), .Y(n1855) );
  NAND2X1 U1822 ( .A(\mem<1><10> ), .B(n159), .Y(n1809) );
  OAI21X1 U1823 ( .A(n158), .B(n1283), .C(n1809), .Y(n1854) );
  NAND2X1 U1824 ( .A(\mem<1><11> ), .B(n159), .Y(n1810) );
  OAI21X1 U1825 ( .A(n158), .B(n1284), .C(n1810), .Y(n1853) );
  NAND2X1 U1826 ( .A(\mem<1><12> ), .B(n159), .Y(n1811) );
  OAI21X1 U1827 ( .A(n158), .B(n1286), .C(n1811), .Y(n1852) );
  NAND2X1 U1828 ( .A(\mem<1><13> ), .B(n159), .Y(n1812) );
  OAI21X1 U1829 ( .A(n158), .B(n1288), .C(n1812), .Y(n1851) );
  NAND2X1 U1830 ( .A(\mem<1><14> ), .B(n159), .Y(n1813) );
  OAI21X1 U1831 ( .A(n158), .B(n1290), .C(n1813), .Y(n1850) );
  NAND2X1 U1832 ( .A(\mem<1><15> ), .B(n159), .Y(n1814) );
  OAI21X1 U1833 ( .A(n158), .B(n1292), .C(n1814), .Y(n1849) );
  NAND2X1 U1834 ( .A(\mem<0><0> ), .B(n1264), .Y(n1817) );
  OAI21X1 U1835 ( .A(n1263), .B(n1270), .C(n1817), .Y(n1848) );
  NAND2X1 U1836 ( .A(\mem<0><1> ), .B(n1264), .Y(n1818) );
  OAI21X1 U1837 ( .A(n1263), .B(n1271), .C(n1818), .Y(n1847) );
  NAND2X1 U1838 ( .A(\mem<0><2> ), .B(n1264), .Y(n1819) );
  OAI21X1 U1839 ( .A(n1263), .B(n1273), .C(n1819), .Y(n1846) );
  NAND2X1 U1840 ( .A(\mem<0><3> ), .B(n1264), .Y(n1820) );
  OAI21X1 U1841 ( .A(n1263), .B(n1274), .C(n1820), .Y(n1845) );
  NAND2X1 U1842 ( .A(\mem<0><4> ), .B(n1264), .Y(n1821) );
  OAI21X1 U1843 ( .A(n1263), .B(n1275), .C(n1821), .Y(n1844) );
  NAND2X1 U1844 ( .A(\mem<0><5> ), .B(n1264), .Y(n1822) );
  OAI21X1 U1845 ( .A(n1263), .B(n1276), .C(n1822), .Y(n1843) );
  NAND2X1 U1846 ( .A(\mem<0><6> ), .B(n1264), .Y(n1823) );
  OAI21X1 U1847 ( .A(n1263), .B(n1278), .C(n1823), .Y(n1842) );
  NAND2X1 U1848 ( .A(\mem<0><7> ), .B(n1264), .Y(n1824) );
  OAI21X1 U1849 ( .A(n1263), .B(n1279), .C(n1824), .Y(n1841) );
  NAND2X1 U1850 ( .A(\mem<0><8> ), .B(n1265), .Y(n1825) );
  OAI21X1 U1851 ( .A(n1263), .B(n1280), .C(n1825), .Y(n1840) );
  NAND2X1 U1852 ( .A(\mem<0><9> ), .B(n1265), .Y(n1826) );
  OAI21X1 U1853 ( .A(n1263), .B(n1281), .C(n1826), .Y(n1839) );
  NAND2X1 U1854 ( .A(\mem<0><10> ), .B(n1265), .Y(n1827) );
  OAI21X1 U1855 ( .A(n1263), .B(n1283), .C(n1827), .Y(n1838) );
  NAND2X1 U1856 ( .A(\mem<0><11> ), .B(n1265), .Y(n1828) );
  OAI21X1 U1857 ( .A(n1263), .B(n1284), .C(n1828), .Y(n1837) );
  NAND2X1 U1858 ( .A(\mem<0><12> ), .B(n1265), .Y(n1829) );
  OAI21X1 U1859 ( .A(n1263), .B(n1286), .C(n1829), .Y(n1836) );
  NAND2X1 U1860 ( .A(\mem<0><13> ), .B(n1265), .Y(n1830) );
  OAI21X1 U1861 ( .A(n1263), .B(n1288), .C(n1830), .Y(n1835) );
  NAND2X1 U1862 ( .A(\mem<0><14> ), .B(n1265), .Y(n1831) );
  OAI21X1 U1863 ( .A(n1263), .B(n1290), .C(n1831), .Y(n1834) );
  NAND2X1 U1864 ( .A(\mem<0><15> ), .B(n1265), .Y(n1832) );
  OAI21X1 U1865 ( .A(n1263), .B(n1292), .C(n1832), .Y(n1833) );
endmodule


module memc_Size16_1 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n1788), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n1789), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n1790), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n1791), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n1792), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n1793), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n1794), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n1795), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n1796), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1797), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1798), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1799), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1800), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1801), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1802), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1803), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n1804), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n1805), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n1806), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n1807), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n1808), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n1809), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n1810), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n1811), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1812), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1813), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1814), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1815), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1816), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1817), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1818), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1819), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n1820), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n1821), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n1822), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n1823), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n1824), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n1825), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n1826), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n1827), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1828), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1829), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1830), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1831), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1832), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1833), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1834), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1835), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n1836), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n1837), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n1838), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n1839), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n1840), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n1841), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n1842), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n1843), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1844), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1845), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1846), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1847), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1848), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1849), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1850), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1851), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n1852), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n1853), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n1854), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n1855), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n1856), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n1857), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n1858), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n1859), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1860), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1861), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1862), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1863), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1864), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1865), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1866), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1867), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n1868), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n1869), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n1870), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n1871), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n1872), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n1873), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n1874), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n1875), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1876), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1877), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1878), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1879), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1880), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1881), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1882), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1883), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n1884), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n1885), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n1886), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n1887), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n1888), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n1889), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n1890), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n1891), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1892), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1893), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1894), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1895), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1896), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1897), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1898), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1899), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n1900), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n1901), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n1902), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n1903), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n1904), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n1905), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n1906), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n1907), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1908), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1909), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1910), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1911), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1912), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1913), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1914), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1915), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n1916), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n1917), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n1918), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n1919), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n1920), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n1921), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n1922), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n1923), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1924), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1925), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1926), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1927), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1928), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1929), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1930), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1931), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n1932), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n1933), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n1934), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n1935), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n1936), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n1937), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n1938), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n1939), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n1940), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n1941), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n1942), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n1943), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n1944), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n1945), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n1946), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n1947), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n1948), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n1949), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n1950), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n1951), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n1952), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n1953), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n1954), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n1955), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n1956), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n1957), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n1958), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n1959), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n1960), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n1961), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n1962), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n1963), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n1964), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n1965), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n1966), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n1967), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n1968), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n1969), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n1970), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n1971), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n1972), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n1973), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n1974), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n1975), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n1976), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n1977), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n1978), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n1979), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n1980), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n1981), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n1982), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n1983), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n1984), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n1985), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n1986), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n1987), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n1988), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n1989), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n1990), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n1991), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n1992), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n1993), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n1994), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n1995), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n1996), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n1997), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n1998), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n1999), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n2000), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n2001), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n2002), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n2003), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2004), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2005), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2006), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2007), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2008), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2009), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2010), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2011), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n2012), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n2013), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n2014), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n2015), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n2016), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n2017), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n2018), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n2019), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2020), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2021), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2022), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2023), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2024), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2025), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2026), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2027), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n2028), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n2029), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n2030), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n2031), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n2032), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n2033), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n2034), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n2035), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2036), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2037), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2038), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2039), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2040), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2041), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2042), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2043), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n2044), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n2045), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n2046), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n2047), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n2048), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n2049), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n2050), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n2051), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2052), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2053), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2054), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2055), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2056), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2057), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2058), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2059), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n2060), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n2061), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n2062), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n2063), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n2064), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n2065), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n2066), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n2067), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2068), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2069), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2070), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2071), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2072), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2073), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2074), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2075), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n2076), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n2077), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n2078), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n2079), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n2080), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n2081), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n2082), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n2083), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2084), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2085), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2086), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2087), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2088), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2089), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2090), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2091), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n2092), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n2093), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n2094), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n2095), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n2096), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n2097), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n2098), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n2099), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2100), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2101), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2102), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2103), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2104), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2105), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2106), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2107), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n2108), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n2109), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n2110), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n2111), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n2112), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n2113), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n2114), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n2115), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2116), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2117), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2118), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2119), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2120), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2121), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2122), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2123), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n2124), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n2125), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n2126), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n2127), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n2128), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n2129), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n2130), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n2131), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2132), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2133), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2134), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2135), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2136), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2137), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2138), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2139), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n2140), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n2141), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n2142), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n2143), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n2144), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n2145), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n2146), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n2147), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2148), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2149), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2150), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2151), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2152), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2153), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2154), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2155), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n2156), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n2157), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n2158), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n2159), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n2160), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n2161), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n2162), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n2163), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2164), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2165), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2166), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2167), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2168), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2169), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2170), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2171), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n2172), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n2173), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n2174), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n2175), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n2176), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n2177), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n2178), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n2179), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2180), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2181), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2182), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2183), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2184), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2185), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2186), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2187), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n2188), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n2189), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n2190), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n2191), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n2192), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n2193), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n2194), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n2195), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2196), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2197), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2198), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2199), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2200), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2201), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2202), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2203), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n2204), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n2205), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n2206), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n2207), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n2208), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n2209), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n2210), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n2211), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2212), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2213), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2214), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2215), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2216), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2217), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2218), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2219), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n2220), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n2221), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n2222), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n2223), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n2224), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n2225), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n2226), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n2227), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2228), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2229), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2230), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2231), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2232), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2233), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2234), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2235), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n2236), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n2237), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n2238), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n2239), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n2240), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n2241), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n2242), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n2243), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2244), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2245), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2246), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2247), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2248), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2249), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2250), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2251), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n2252), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n2253), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n2254), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n2255), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n2256), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n2257), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n2258), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n2259), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2260), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2261), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2262), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2263), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2264), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2265), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2266), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2267), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n2268), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n2269), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n2270), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n2271), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n2272), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n2273), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n2274), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n2275), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2276), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2277), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2278), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2279), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2280), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2281), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2282), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2283), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n2284), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n2285), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n2286), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n2287), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n2288), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n2289), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n2290), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n2291), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2292), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2293), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2294), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2295), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2296), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2297), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2298), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2299), .CLK(clk), .Q(\mem<31><0> ) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n2300) );
  INVX4 U2 ( .A(n27), .Y(n136) );
  INVX1 U3 ( .A(n1207), .Y(n1192) );
  INVX1 U4 ( .A(n1191), .Y(n1201) );
  INVX1 U5 ( .A(n1191), .Y(n1200) );
  INVX1 U6 ( .A(n1191), .Y(n1202) );
  INVX1 U7 ( .A(n1191), .Y(n1203) );
  INVX1 U8 ( .A(n1192), .Y(n1199) );
  INVX1 U9 ( .A(n1191), .Y(n1205) );
  INVX1 U10 ( .A(n1192), .Y(n1197) );
  INVX1 U11 ( .A(n1192), .Y(n1196) );
  AND2X2 U12 ( .A(n1251), .B(n48), .Y(n59) );
  INVX1 U13 ( .A(n640), .Y(N32) );
  INVX1 U14 ( .A(n641), .Y(N31) );
  INVX1 U15 ( .A(n642), .Y(N30) );
  INVX1 U16 ( .A(n643), .Y(N29) );
  INVX1 U17 ( .A(n644), .Y(N28) );
  INVX1 U18 ( .A(n645), .Y(N27) );
  INVX1 U19 ( .A(n646), .Y(N26) );
  INVX1 U20 ( .A(n647), .Y(N25) );
  INVX1 U21 ( .A(n648), .Y(N24) );
  INVX1 U22 ( .A(n650), .Y(N22) );
  INVX1 U23 ( .A(n1163), .Y(N21) );
  INVX1 U24 ( .A(n1165), .Y(N19) );
  INVX1 U25 ( .A(n1166), .Y(N18) );
  INVX1 U26 ( .A(n1167), .Y(N17) );
  INVX1 U27 ( .A(n1251), .Y(n1207) );
  INVX1 U28 ( .A(N10), .Y(n1191) );
  INVX1 U29 ( .A(n1192), .Y(n1193) );
  INVX1 U30 ( .A(n1190), .Y(n1179) );
  INVX2 U31 ( .A(n1191), .Y(n1194) );
  INVX1 U32 ( .A(n1190), .Y(n1180) );
  INVX1 U33 ( .A(n1171), .Y(n1176) );
  INVX2 U34 ( .A(n1191), .Y(n1195) );
  INVX1 U35 ( .A(n1190), .Y(n1181) );
  INVX1 U36 ( .A(n1178), .Y(n1182) );
  INVX2 U37 ( .A(n1192), .Y(n1198) );
  INVX1 U38 ( .A(n1178), .Y(n1183) );
  INVX1 U39 ( .A(n1178), .Y(n1184) );
  INVX1 U40 ( .A(n1171), .Y(n1174) );
  INVX1 U41 ( .A(n1177), .Y(n1185) );
  INVX1 U42 ( .A(n1177), .Y(n1186) );
  INVX2 U43 ( .A(n1191), .Y(n1204) );
  INVX1 U44 ( .A(n1177), .Y(n1187) );
  INVX1 U45 ( .A(n1178), .Y(n1188) );
  INVX2 U46 ( .A(n1251), .Y(n1206) );
  INVX1 U47 ( .A(n1177), .Y(n1189) );
  INVX1 U48 ( .A(n649), .Y(N23) );
  INVX1 U49 ( .A(n1164), .Y(N20) );
  INVX1 U50 ( .A(n1252), .Y(n1190) );
  INVX1 U51 ( .A(n1254), .Y(n1171) );
  INVX1 U52 ( .A(n1171), .Y(n1173) );
  INVX1 U53 ( .A(n1171), .Y(n1175) );
  INVX1 U54 ( .A(n1171), .Y(n1172) );
  INVX1 U55 ( .A(N14), .Y(n1258) );
  INVX1 U56 ( .A(n1256), .Y(n1169) );
  INVX1 U57 ( .A(n1256), .Y(n1170) );
  INVX1 U58 ( .A(n1258), .Y(n1168) );
  INVX1 U59 ( .A(rst), .Y(n1249) );
  INVX1 U60 ( .A(n1252), .Y(n1177) );
  INVX1 U61 ( .A(n1252), .Y(n1178) );
  INVX1 U62 ( .A(n66), .Y(n1208) );
  INVX1 U63 ( .A(n67), .Y(n1209) );
  INVX1 U64 ( .A(n68), .Y(n1210) );
  INVX4 U65 ( .A(n4), .Y(n73) );
  INVX4 U66 ( .A(n15), .Y(n104) );
  INVX4 U67 ( .A(n14), .Y(n101) );
  INVX4 U68 ( .A(n13), .Y(n98) );
  INVX4 U69 ( .A(n12), .Y(n95) );
  INVX4 U70 ( .A(n10), .Y(n91) );
  INVX4 U71 ( .A(n9), .Y(n88) );
  INVX4 U72 ( .A(n8), .Y(n85) );
  INVX4 U73 ( .A(n7), .Y(n82) );
  INVX4 U74 ( .A(n6), .Y(n79) );
  INVX4 U75 ( .A(n5), .Y(n76) );
  INVX4 U76 ( .A(n11), .Y(n92) );
  INVX4 U77 ( .A(n1215), .Y(n1214) );
  INVX4 U78 ( .A(n26), .Y(n135) );
  INVX4 U79 ( .A(n25), .Y(n132) );
  INVX4 U80 ( .A(n24), .Y(n129) );
  INVX4 U81 ( .A(n23), .Y(n126) );
  INVX4 U82 ( .A(n22), .Y(n123) );
  INVX4 U83 ( .A(n21), .Y(n120) );
  INVX4 U84 ( .A(n20), .Y(n117) );
  INVX4 U85 ( .A(n18), .Y(n113) );
  INVX4 U86 ( .A(n17), .Y(n110) );
  INVX4 U87 ( .A(n16), .Y(n107) );
  INVX4 U88 ( .A(n19), .Y(n114) );
  INVX4 U89 ( .A(n35), .Y(n158) );
  INVX4 U90 ( .A(n34), .Y(n157) );
  INVX4 U91 ( .A(n33), .Y(n154) );
  INVX4 U92 ( .A(n32), .Y(n151) );
  INVX4 U93 ( .A(n31), .Y(n148) );
  INVX4 U94 ( .A(n30), .Y(n145) );
  INVX4 U95 ( .A(n29), .Y(n142) );
  INVX4 U96 ( .A(n28), .Y(n139) );
  INVX1 U97 ( .A(n1259), .Y(n1) );
  INVX2 U98 ( .A(n47), .Y(n1216) );
  INVX4 U99 ( .A(n47), .Y(n1215) );
  INVX1 U100 ( .A(n1259), .Y(n1260) );
  BUFX2 U101 ( .A(write), .Y(n2) );
  INVX2 U102 ( .A(n1259), .Y(n3) );
  INVX1 U103 ( .A(N13), .Y(n1256) );
  AND2X2 U104 ( .A(n1211), .B(n71), .Y(n4) );
  AND2X2 U105 ( .A(n1211), .B(n74), .Y(n5) );
  AND2X2 U106 ( .A(n1211), .B(n77), .Y(n6) );
  AND2X2 U107 ( .A(n1211), .B(n80), .Y(n7) );
  AND2X2 U108 ( .A(n1211), .B(n83), .Y(n8) );
  AND2X2 U109 ( .A(n1211), .B(n86), .Y(n9) );
  AND2X2 U110 ( .A(n1211), .B(n89), .Y(n10) );
  AND2X2 U111 ( .A(n1211), .B(n66), .Y(n11) );
  AND2X2 U112 ( .A(n1211), .B(n93), .Y(n12) );
  AND2X2 U113 ( .A(n1211), .B(n96), .Y(n13) );
  AND2X2 U114 ( .A(n1211), .B(n99), .Y(n14) );
  AND2X2 U115 ( .A(n1211), .B(n102), .Y(n15) );
  AND2X2 U116 ( .A(n1212), .B(n105), .Y(n16) );
  AND2X2 U117 ( .A(n1212), .B(n108), .Y(n17) );
  AND2X2 U118 ( .A(n1212), .B(n111), .Y(n18) );
  AND2X2 U119 ( .A(n1212), .B(n67), .Y(n19) );
  AND2X2 U120 ( .A(n1212), .B(n115), .Y(n20) );
  AND2X2 U121 ( .A(n1212), .B(n118), .Y(n21) );
  AND2X2 U122 ( .A(n1212), .B(n121), .Y(n22) );
  AND2X2 U123 ( .A(n1212), .B(n124), .Y(n23) );
  AND2X2 U124 ( .A(n1212), .B(n127), .Y(n24) );
  AND2X2 U125 ( .A(n1212), .B(n130), .Y(n25) );
  AND2X2 U126 ( .A(n1212), .B(n133), .Y(n26) );
  AND2X2 U127 ( .A(n1213), .B(n68), .Y(n27) );
  AND2X2 U128 ( .A(n1213), .B(n137), .Y(n28) );
  AND2X2 U129 ( .A(n1213), .B(n140), .Y(n29) );
  AND2X2 U130 ( .A(n1213), .B(n143), .Y(n30) );
  AND2X2 U131 ( .A(n1213), .B(n146), .Y(n31) );
  AND2X2 U132 ( .A(n1213), .B(n149), .Y(n32) );
  AND2X2 U133 ( .A(n1213), .B(n152), .Y(n33) );
  AND2X2 U134 ( .A(n1213), .B(n155), .Y(n34) );
  AND2X2 U135 ( .A(n1212), .B(n69), .Y(n35) );
  AND2X2 U136 ( .A(\data_in<0> ), .B(n1214), .Y(n36) );
  AND2X2 U137 ( .A(\data_in<1> ), .B(n1214), .Y(n37) );
  AND2X2 U138 ( .A(\data_in<2> ), .B(n1214), .Y(n38) );
  AND2X2 U139 ( .A(\data_in<3> ), .B(n1214), .Y(n39) );
  AND2X2 U140 ( .A(\data_in<4> ), .B(n1214), .Y(n40) );
  AND2X2 U141 ( .A(\data_in<5> ), .B(n1214), .Y(n41) );
  AND2X2 U142 ( .A(\data_in<6> ), .B(n1214), .Y(n42) );
  AND2X2 U143 ( .A(\data_in<7> ), .B(n1214), .Y(n43) );
  AND2X2 U144 ( .A(\data_in<8> ), .B(n1214), .Y(n44) );
  AND2X2 U145 ( .A(\data_in<9> ), .B(n1214), .Y(n45) );
  AND2X2 U146 ( .A(\data_in<10> ), .B(n1214), .Y(n46) );
  AND2X2 U147 ( .A(n2), .B(n1249), .Y(n47) );
  INVX1 U148 ( .A(n1253), .Y(n1252) );
  INVX1 U149 ( .A(n1251), .Y(n1250) );
  AND2X1 U150 ( .A(n1254), .B(n1252), .Y(n48) );
  INVX1 U151 ( .A(n1255), .Y(n1254) );
  AND2X1 U152 ( .A(n2300), .B(n1257), .Y(n49) );
  INVX1 U153 ( .A(n1258), .Y(n1257) );
  BUFX2 U154 ( .A(n1293), .Y(n50) );
  INVX1 U155 ( .A(n50), .Y(n1685) );
  BUFX2 U156 ( .A(n1310), .Y(n51) );
  INVX1 U157 ( .A(n51), .Y(n1702) );
  BUFX2 U158 ( .A(n1327), .Y(n52) );
  INVX1 U159 ( .A(n52), .Y(n1719) );
  BUFX2 U160 ( .A(n1344), .Y(n53) );
  INVX1 U161 ( .A(n53), .Y(n1736) );
  BUFX2 U162 ( .A(n1361), .Y(n54) );
  INVX1 U163 ( .A(n54), .Y(n1753) );
  BUFX2 U164 ( .A(n1522), .Y(n55) );
  INVX1 U165 ( .A(n55), .Y(n1635) );
  BUFX2 U166 ( .A(n1652), .Y(n56) );
  INVX1 U167 ( .A(n56), .Y(n1770) );
  AND2X1 U168 ( .A(n1250), .B(n48), .Y(n57) );
  AND2X1 U169 ( .A(n1170), .B(n49), .Y(n58) );
  AND2X1 U170 ( .A(n1256), .B(n49), .Y(n60) );
  AND2X2 U171 ( .A(\data_in<11> ), .B(n1213), .Y(n61) );
  AND2X2 U172 ( .A(\data_in<12> ), .B(n1213), .Y(n62) );
  AND2X2 U173 ( .A(\data_in<13> ), .B(n1213), .Y(n63) );
  AND2X2 U174 ( .A(\data_in<14> ), .B(n1213), .Y(n64) );
  AND2X2 U175 ( .A(\data_in<15> ), .B(n1213), .Y(n65) );
  AND2X1 U176 ( .A(n58), .B(n1771), .Y(n66) );
  AND2X1 U177 ( .A(n1771), .B(n60), .Y(n67) );
  AND2X1 U178 ( .A(n1771), .B(n1635), .Y(n68) );
  AND2X1 U179 ( .A(n1771), .B(n1770), .Y(n69) );
  INVX1 U180 ( .A(n69), .Y(n70) );
  AND2X1 U181 ( .A(n57), .B(n58), .Y(n71) );
  INVX1 U182 ( .A(n71), .Y(n72) );
  AND2X1 U183 ( .A(n58), .B(n59), .Y(n74) );
  INVX1 U184 ( .A(n74), .Y(n75) );
  AND2X1 U185 ( .A(n58), .B(n1685), .Y(n77) );
  INVX1 U186 ( .A(n77), .Y(n78) );
  AND2X1 U187 ( .A(n58), .B(n1702), .Y(n80) );
  INVX1 U188 ( .A(n80), .Y(n81) );
  AND2X1 U189 ( .A(n58), .B(n1719), .Y(n83) );
  INVX1 U190 ( .A(n83), .Y(n84) );
  AND2X1 U191 ( .A(n58), .B(n1736), .Y(n86) );
  INVX1 U192 ( .A(n86), .Y(n87) );
  AND2X1 U193 ( .A(n58), .B(n1753), .Y(n89) );
  INVX1 U194 ( .A(n89), .Y(n90) );
  AND2X1 U195 ( .A(n57), .B(n60), .Y(n93) );
  INVX1 U196 ( .A(n93), .Y(n94) );
  AND2X1 U197 ( .A(n59), .B(n60), .Y(n96) );
  INVX1 U198 ( .A(n96), .Y(n97) );
  AND2X1 U199 ( .A(n1685), .B(n60), .Y(n99) );
  INVX1 U200 ( .A(n99), .Y(n100) );
  AND2X1 U201 ( .A(n1702), .B(n60), .Y(n102) );
  INVX1 U202 ( .A(n102), .Y(n103) );
  AND2X1 U203 ( .A(n1719), .B(n60), .Y(n105) );
  INVX1 U204 ( .A(n105), .Y(n106) );
  AND2X1 U205 ( .A(n1736), .B(n60), .Y(n108) );
  INVX1 U206 ( .A(n108), .Y(n109) );
  AND2X1 U207 ( .A(n1753), .B(n60), .Y(n111) );
  INVX1 U208 ( .A(n111), .Y(n112) );
  AND2X1 U209 ( .A(n57), .B(n1635), .Y(n115) );
  INVX1 U210 ( .A(n115), .Y(n116) );
  AND2X1 U211 ( .A(n59), .B(n1635), .Y(n118) );
  INVX1 U212 ( .A(n118), .Y(n119) );
  AND2X1 U213 ( .A(n1685), .B(n1635), .Y(n121) );
  INVX1 U214 ( .A(n121), .Y(n122) );
  AND2X1 U215 ( .A(n1702), .B(n1635), .Y(n124) );
  INVX1 U216 ( .A(n124), .Y(n125) );
  AND2X1 U217 ( .A(n1719), .B(n1635), .Y(n127) );
  INVX1 U218 ( .A(n127), .Y(n128) );
  AND2X1 U219 ( .A(n1736), .B(n1635), .Y(n130) );
  INVX1 U220 ( .A(n130), .Y(n131) );
  AND2X1 U221 ( .A(n1753), .B(n1635), .Y(n133) );
  INVX1 U222 ( .A(n133), .Y(n134) );
  AND2X1 U223 ( .A(n57), .B(n1770), .Y(n137) );
  INVX1 U224 ( .A(n137), .Y(n138) );
  AND2X1 U225 ( .A(n59), .B(n1770), .Y(n140) );
  INVX1 U226 ( .A(n140), .Y(n141) );
  AND2X1 U227 ( .A(n1685), .B(n1770), .Y(n143) );
  INVX1 U228 ( .A(n143), .Y(n144) );
  AND2X1 U229 ( .A(n1702), .B(n1770), .Y(n146) );
  INVX1 U230 ( .A(n146), .Y(n147) );
  AND2X1 U231 ( .A(n1719), .B(n1770), .Y(n149) );
  INVX1 U232 ( .A(n149), .Y(n150) );
  AND2X1 U233 ( .A(n1736), .B(n1770), .Y(n152) );
  INVX1 U234 ( .A(n152), .Y(n153) );
  AND2X1 U235 ( .A(n1753), .B(n1770), .Y(n155) );
  INVX1 U236 ( .A(n155), .Y(n156) );
  MUX2X1 U237 ( .B(n160), .A(n161), .S(n1179), .Y(n159) );
  MUX2X1 U238 ( .B(n163), .A(n164), .S(n1179), .Y(n162) );
  MUX2X1 U239 ( .B(n166), .A(n167), .S(n1179), .Y(n165) );
  MUX2X1 U240 ( .B(n169), .A(n170), .S(n1179), .Y(n168) );
  MUX2X1 U241 ( .B(n172), .A(n173), .S(n1170), .Y(n171) );
  MUX2X1 U242 ( .B(n175), .A(n176), .S(n1179), .Y(n174) );
  MUX2X1 U243 ( .B(n178), .A(n179), .S(n1179), .Y(n177) );
  MUX2X1 U244 ( .B(n181), .A(n182), .S(n1179), .Y(n180) );
  MUX2X1 U245 ( .B(n184), .A(n185), .S(n1179), .Y(n183) );
  MUX2X1 U246 ( .B(n187), .A(n188), .S(n1170), .Y(n186) );
  MUX2X1 U247 ( .B(n190), .A(n191), .S(n1180), .Y(n189) );
  MUX2X1 U248 ( .B(n193), .A(n194), .S(n1180), .Y(n192) );
  MUX2X1 U249 ( .B(n196), .A(n197), .S(n1180), .Y(n195) );
  MUX2X1 U250 ( .B(n199), .A(n200), .S(n1180), .Y(n198) );
  MUX2X1 U251 ( .B(n202), .A(n203), .S(n1170), .Y(n201) );
  MUX2X1 U252 ( .B(n205), .A(n206), .S(n1180), .Y(n204) );
  MUX2X1 U253 ( .B(n208), .A(n209), .S(n1180), .Y(n207) );
  MUX2X1 U254 ( .B(n211), .A(n212), .S(n1180), .Y(n210) );
  MUX2X1 U255 ( .B(n215), .A(n216), .S(n1180), .Y(n213) );
  MUX2X1 U256 ( .B(n218), .A(n219), .S(n1170), .Y(n217) );
  MUX2X1 U257 ( .B(n221), .A(n222), .S(n1180), .Y(n220) );
  MUX2X1 U258 ( .B(n224), .A(n225), .S(n1180), .Y(n223) );
  MUX2X1 U259 ( .B(n227), .A(n228), .S(n1180), .Y(n226) );
  MUX2X1 U260 ( .B(n230), .A(n231), .S(n1180), .Y(n229) );
  MUX2X1 U261 ( .B(n233), .A(n234), .S(n1170), .Y(n232) );
  MUX2X1 U262 ( .B(n236), .A(n237), .S(n1181), .Y(n235) );
  MUX2X1 U263 ( .B(n239), .A(n240), .S(n1181), .Y(n238) );
  MUX2X1 U264 ( .B(n242), .A(n243), .S(n1181), .Y(n241) );
  MUX2X1 U265 ( .B(n245), .A(n246), .S(n1181), .Y(n244) );
  MUX2X1 U266 ( .B(n248), .A(n249), .S(n1170), .Y(n247) );
  MUX2X1 U267 ( .B(n251), .A(n252), .S(n1181), .Y(n250) );
  MUX2X1 U268 ( .B(n254), .A(n255), .S(n1181), .Y(n253) );
  MUX2X1 U269 ( .B(n257), .A(n258), .S(n1181), .Y(n256) );
  MUX2X1 U270 ( .B(n260), .A(n261), .S(n1181), .Y(n259) );
  MUX2X1 U271 ( .B(n263), .A(n264), .S(n1170), .Y(n262) );
  MUX2X1 U272 ( .B(n266), .A(n267), .S(n1181), .Y(n265) );
  MUX2X1 U273 ( .B(n269), .A(n270), .S(n1181), .Y(n268) );
  MUX2X1 U274 ( .B(n272), .A(n273), .S(n1181), .Y(n271) );
  MUX2X1 U275 ( .B(n275), .A(n276), .S(n1181), .Y(n274) );
  MUX2X1 U276 ( .B(n278), .A(n279), .S(n1170), .Y(n277) );
  MUX2X1 U277 ( .B(n281), .A(n282), .S(n1182), .Y(n280) );
  MUX2X1 U278 ( .B(n284), .A(n285), .S(n1182), .Y(n283) );
  MUX2X1 U279 ( .B(n287), .A(n288), .S(n1182), .Y(n286) );
  MUX2X1 U280 ( .B(n290), .A(n291), .S(n1182), .Y(n289) );
  MUX2X1 U281 ( .B(n293), .A(n294), .S(n1170), .Y(n292) );
  MUX2X1 U282 ( .B(n296), .A(n297), .S(n1182), .Y(n295) );
  MUX2X1 U283 ( .B(n299), .A(n300), .S(n1182), .Y(n298) );
  MUX2X1 U284 ( .B(n302), .A(n303), .S(n1182), .Y(n301) );
  MUX2X1 U285 ( .B(n305), .A(n306), .S(n1182), .Y(n304) );
  MUX2X1 U286 ( .B(n308), .A(n309), .S(n1170), .Y(n307) );
  MUX2X1 U287 ( .B(n311), .A(n312), .S(n1182), .Y(n310) );
  MUX2X1 U288 ( .B(n314), .A(n315), .S(n1182), .Y(n313) );
  MUX2X1 U289 ( .B(n317), .A(n318), .S(n1182), .Y(n316) );
  MUX2X1 U290 ( .B(n320), .A(n321), .S(n1182), .Y(n319) );
  MUX2X1 U291 ( .B(n323), .A(n324), .S(n1170), .Y(n322) );
  MUX2X1 U292 ( .B(n326), .A(n327), .S(n1183), .Y(n325) );
  MUX2X1 U293 ( .B(n329), .A(n330), .S(n1183), .Y(n328) );
  MUX2X1 U294 ( .B(n332), .A(n333), .S(n1183), .Y(n331) );
  MUX2X1 U295 ( .B(n335), .A(n336), .S(n1183), .Y(n334) );
  MUX2X1 U296 ( .B(n338), .A(n339), .S(n1170), .Y(n337) );
  MUX2X1 U297 ( .B(n341), .A(n342), .S(n1183), .Y(n340) );
  MUX2X1 U298 ( .B(n344), .A(n345), .S(n1183), .Y(n343) );
  MUX2X1 U299 ( .B(n347), .A(n348), .S(n1183), .Y(n346) );
  MUX2X1 U300 ( .B(n350), .A(n351), .S(n1183), .Y(n349) );
  MUX2X1 U301 ( .B(n353), .A(n354), .S(n1169), .Y(n352) );
  MUX2X1 U302 ( .B(n356), .A(n357), .S(n1183), .Y(n355) );
  MUX2X1 U303 ( .B(n359), .A(n360), .S(n1183), .Y(n358) );
  MUX2X1 U304 ( .B(n362), .A(n363), .S(n1183), .Y(n361) );
  MUX2X1 U305 ( .B(n365), .A(n366), .S(n1183), .Y(n364) );
  MUX2X1 U306 ( .B(n368), .A(n369), .S(n1169), .Y(n367) );
  MUX2X1 U307 ( .B(n371), .A(n372), .S(n1184), .Y(n370) );
  MUX2X1 U308 ( .B(n374), .A(n375), .S(n1184), .Y(n373) );
  MUX2X1 U309 ( .B(n377), .A(n378), .S(n1184), .Y(n376) );
  MUX2X1 U310 ( .B(n380), .A(n381), .S(n1184), .Y(n379) );
  MUX2X1 U311 ( .B(n383), .A(n384), .S(n1169), .Y(n382) );
  MUX2X1 U312 ( .B(n386), .A(n387), .S(n1184), .Y(n385) );
  MUX2X1 U313 ( .B(n389), .A(n390), .S(n1184), .Y(n388) );
  MUX2X1 U314 ( .B(n392), .A(n393), .S(n1184), .Y(n391) );
  MUX2X1 U315 ( .B(n395), .A(n396), .S(n1184), .Y(n394) );
  MUX2X1 U316 ( .B(n398), .A(n399), .S(n1169), .Y(n397) );
  MUX2X1 U317 ( .B(n401), .A(n402), .S(n1184), .Y(n400) );
  MUX2X1 U318 ( .B(n404), .A(n405), .S(n1184), .Y(n403) );
  MUX2X1 U319 ( .B(n407), .A(n408), .S(n1184), .Y(n406) );
  MUX2X1 U320 ( .B(n410), .A(n411), .S(n1184), .Y(n409) );
  MUX2X1 U321 ( .B(n413), .A(n414), .S(n1169), .Y(n412) );
  MUX2X1 U322 ( .B(n416), .A(n417), .S(n1185), .Y(n415) );
  MUX2X1 U323 ( .B(n419), .A(n420), .S(n1185), .Y(n418) );
  MUX2X1 U324 ( .B(n422), .A(n423), .S(n1185), .Y(n421) );
  MUX2X1 U325 ( .B(n425), .A(n426), .S(n1185), .Y(n424) );
  MUX2X1 U326 ( .B(n428), .A(n429), .S(n1169), .Y(n427) );
  MUX2X1 U327 ( .B(n431), .A(n432), .S(n1185), .Y(n430) );
  MUX2X1 U328 ( .B(n434), .A(n435), .S(n1185), .Y(n433) );
  MUX2X1 U329 ( .B(n437), .A(n438), .S(n1185), .Y(n436) );
  MUX2X1 U330 ( .B(n440), .A(n441), .S(n1185), .Y(n439) );
  MUX2X1 U331 ( .B(n443), .A(n444), .S(n1169), .Y(n442) );
  MUX2X1 U332 ( .B(n446), .A(n447), .S(n1185), .Y(n445) );
  MUX2X1 U333 ( .B(n449), .A(n450), .S(n1185), .Y(n448) );
  MUX2X1 U334 ( .B(n452), .A(n453), .S(n1185), .Y(n451) );
  MUX2X1 U335 ( .B(n455), .A(n456), .S(n1185), .Y(n454) );
  MUX2X1 U336 ( .B(n458), .A(n459), .S(n1169), .Y(n457) );
  MUX2X1 U337 ( .B(n461), .A(n462), .S(n1186), .Y(n460) );
  MUX2X1 U338 ( .B(n464), .A(n465), .S(n1186), .Y(n463) );
  MUX2X1 U339 ( .B(n467), .A(n468), .S(n1186), .Y(n466) );
  MUX2X1 U340 ( .B(n470), .A(n471), .S(n1186), .Y(n469) );
  MUX2X1 U341 ( .B(n473), .A(n474), .S(n1169), .Y(n472) );
  MUX2X1 U342 ( .B(n476), .A(n477), .S(n1186), .Y(n475) );
  MUX2X1 U343 ( .B(n479), .A(n480), .S(n1186), .Y(n478) );
  MUX2X1 U344 ( .B(n482), .A(n483), .S(n1186), .Y(n481) );
  MUX2X1 U345 ( .B(n485), .A(n486), .S(n1186), .Y(n484) );
  MUX2X1 U346 ( .B(n488), .A(n489), .S(n1169), .Y(n487) );
  MUX2X1 U347 ( .B(n491), .A(n492), .S(n1186), .Y(n490) );
  MUX2X1 U348 ( .B(n494), .A(n495), .S(n1186), .Y(n493) );
  MUX2X1 U349 ( .B(n497), .A(n498), .S(n1186), .Y(n496) );
  MUX2X1 U350 ( .B(n500), .A(n501), .S(n1186), .Y(n499) );
  MUX2X1 U351 ( .B(n503), .A(n504), .S(n1169), .Y(n502) );
  MUX2X1 U352 ( .B(n506), .A(n507), .S(n1187), .Y(n505) );
  MUX2X1 U353 ( .B(n509), .A(n510), .S(n1187), .Y(n508) );
  MUX2X1 U354 ( .B(n512), .A(n513), .S(n1187), .Y(n511) );
  MUX2X1 U355 ( .B(n515), .A(n516), .S(n1187), .Y(n514) );
  MUX2X1 U356 ( .B(n518), .A(n519), .S(n1169), .Y(n517) );
  MUX2X1 U357 ( .B(n521), .A(n522), .S(n1187), .Y(n520) );
  MUX2X1 U358 ( .B(n524), .A(n525), .S(n1187), .Y(n523) );
  MUX2X1 U359 ( .B(n527), .A(n528), .S(n1187), .Y(n526) );
  MUX2X1 U360 ( .B(n530), .A(n531), .S(n1187), .Y(n529) );
  MUX2X1 U361 ( .B(n533), .A(n534), .S(n1169), .Y(n532) );
  MUX2X1 U362 ( .B(n536), .A(n537), .S(n1187), .Y(n535) );
  MUX2X1 U363 ( .B(n539), .A(n540), .S(n1187), .Y(n538) );
  MUX2X1 U364 ( .B(n542), .A(n543), .S(n1187), .Y(n541) );
  MUX2X1 U365 ( .B(n545), .A(n546), .S(n1187), .Y(n544) );
  MUX2X1 U366 ( .B(n548), .A(n549), .S(n1169), .Y(n547) );
  MUX2X1 U367 ( .B(n551), .A(n552), .S(n1188), .Y(n550) );
  MUX2X1 U368 ( .B(n554), .A(n555), .S(n1188), .Y(n553) );
  MUX2X1 U369 ( .B(n557), .A(n558), .S(n1188), .Y(n556) );
  MUX2X1 U370 ( .B(n560), .A(n561), .S(n1188), .Y(n559) );
  MUX2X1 U371 ( .B(n563), .A(n564), .S(n1169), .Y(n562) );
  MUX2X1 U372 ( .B(n566), .A(n567), .S(n1188), .Y(n565) );
  MUX2X1 U373 ( .B(n569), .A(n570), .S(n1188), .Y(n568) );
  MUX2X1 U374 ( .B(n572), .A(n573), .S(n1188), .Y(n571) );
  MUX2X1 U375 ( .B(n575), .A(n576), .S(n1188), .Y(n574) );
  MUX2X1 U376 ( .B(n578), .A(n579), .S(n1169), .Y(n577) );
  MUX2X1 U377 ( .B(n581), .A(n582), .S(n1188), .Y(n580) );
  MUX2X1 U378 ( .B(n584), .A(n585), .S(n1188), .Y(n583) );
  MUX2X1 U379 ( .B(n587), .A(n588), .S(n1188), .Y(n586) );
  MUX2X1 U380 ( .B(n590), .A(n591), .S(n1188), .Y(n589) );
  MUX2X1 U381 ( .B(n593), .A(n594), .S(n1169), .Y(n592) );
  MUX2X1 U382 ( .B(n596), .A(n597), .S(n1189), .Y(n595) );
  MUX2X1 U383 ( .B(n599), .A(n600), .S(n1189), .Y(n598) );
  MUX2X1 U384 ( .B(n602), .A(n603), .S(n1189), .Y(n601) );
  MUX2X1 U385 ( .B(n605), .A(n606), .S(n1189), .Y(n604) );
  MUX2X1 U386 ( .B(n608), .A(n609), .S(n1169), .Y(n607) );
  MUX2X1 U387 ( .B(n611), .A(n612), .S(n1189), .Y(n610) );
  MUX2X1 U388 ( .B(n614), .A(n615), .S(n1189), .Y(n613) );
  MUX2X1 U389 ( .B(n617), .A(n618), .S(n1189), .Y(n616) );
  MUX2X1 U390 ( .B(n620), .A(n621), .S(n1189), .Y(n619) );
  MUX2X1 U391 ( .B(n623), .A(n624), .S(n1170), .Y(n622) );
  MUX2X1 U392 ( .B(n626), .A(n627), .S(n1189), .Y(n625) );
  MUX2X1 U393 ( .B(n629), .A(n630), .S(n1189), .Y(n628) );
  MUX2X1 U394 ( .B(n632), .A(n633), .S(n1189), .Y(n631) );
  MUX2X1 U395 ( .B(n635), .A(n636), .S(n1189), .Y(n634) );
  MUX2X1 U396 ( .B(n638), .A(n639), .S(n1169), .Y(n637) );
  MUX2X1 U397 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n1193), .Y(n161) );
  MUX2X1 U398 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n1193), .Y(n160) );
  MUX2X1 U399 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n1193), .Y(n164) );
  MUX2X1 U400 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n1193), .Y(n163) );
  MUX2X1 U401 ( .B(n162), .A(n159), .S(n1176), .Y(n173) );
  MUX2X1 U402 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n1196), .Y(n167) );
  MUX2X1 U403 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n1197), .Y(n166) );
  MUX2X1 U404 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n1250), .Y(n170) );
  MUX2X1 U405 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n1205), .Y(n169) );
  MUX2X1 U406 ( .B(n168), .A(n165), .S(n1176), .Y(n172) );
  MUX2X1 U407 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n1250), .Y(n176) );
  MUX2X1 U408 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n1195), .Y(n175) );
  MUX2X1 U409 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n1250), .Y(n179) );
  MUX2X1 U410 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n1250), .Y(n178) );
  MUX2X1 U411 ( .B(n177), .A(n174), .S(n1176), .Y(n188) );
  MUX2X1 U412 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n1194), .Y(n182) );
  MUX2X1 U413 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n1193), .Y(n181) );
  MUX2X1 U414 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n1250), .Y(n185) );
  MUX2X1 U415 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n1250), .Y(n184) );
  MUX2X1 U416 ( .B(n183), .A(n180), .S(n1176), .Y(n187) );
  MUX2X1 U417 ( .B(n186), .A(n171), .S(n1168), .Y(n640) );
  MUX2X1 U418 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n1194), .Y(n191) );
  MUX2X1 U419 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n1194), .Y(n190) );
  MUX2X1 U420 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n1194), .Y(n194) );
  MUX2X1 U421 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n1194), .Y(n193) );
  MUX2X1 U422 ( .B(n192), .A(n189), .S(n1176), .Y(n203) );
  MUX2X1 U423 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n1194), .Y(n197) );
  MUX2X1 U424 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n1194), .Y(n196) );
  MUX2X1 U425 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n1194), .Y(n200) );
  MUX2X1 U426 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n1194), .Y(n199) );
  MUX2X1 U427 ( .B(n198), .A(n195), .S(n1176), .Y(n202) );
  MUX2X1 U428 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n1194), .Y(n206) );
  MUX2X1 U429 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n1194), .Y(n205) );
  MUX2X1 U430 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n1194), .Y(n209) );
  MUX2X1 U431 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n1194), .Y(n208) );
  MUX2X1 U432 ( .B(n207), .A(n204), .S(n1176), .Y(n219) );
  MUX2X1 U433 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n1203), .Y(n212) );
  MUX2X1 U434 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n1250), .Y(n211) );
  MUX2X1 U435 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n1195), .Y(n216) );
  MUX2X1 U436 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n1250), .Y(n215) );
  MUX2X1 U437 ( .B(n213), .A(n210), .S(n1176), .Y(n218) );
  MUX2X1 U438 ( .B(n217), .A(n201), .S(n1168), .Y(n641) );
  MUX2X1 U439 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n1204), .Y(n222) );
  MUX2X1 U440 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n1205), .Y(n221) );
  MUX2X1 U441 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n1204), .Y(n225) );
  MUX2X1 U442 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n1195), .Y(n224) );
  MUX2X1 U443 ( .B(n223), .A(n220), .S(n1176), .Y(n234) );
  MUX2X1 U444 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n1199), .Y(n228) );
  MUX2X1 U445 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n1203), .Y(n227) );
  MUX2X1 U446 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n1195), .Y(n231) );
  MUX2X1 U447 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n1204), .Y(n230) );
  MUX2X1 U448 ( .B(n229), .A(n226), .S(n1176), .Y(n233) );
  MUX2X1 U449 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n1195), .Y(n237) );
  MUX2X1 U450 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n1195), .Y(n236) );
  MUX2X1 U451 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n1195), .Y(n240) );
  MUX2X1 U452 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n1195), .Y(n239) );
  MUX2X1 U453 ( .B(n238), .A(n235), .S(n1176), .Y(n249) );
  MUX2X1 U454 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n1195), .Y(n243) );
  MUX2X1 U455 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n1195), .Y(n242) );
  MUX2X1 U456 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n1195), .Y(n246) );
  MUX2X1 U457 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n1195), .Y(n245) );
  MUX2X1 U458 ( .B(n244), .A(n241), .S(n1176), .Y(n248) );
  MUX2X1 U459 ( .B(n247), .A(n232), .S(n1168), .Y(n642) );
  MUX2X1 U460 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n1195), .Y(n252) );
  MUX2X1 U461 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n1195), .Y(n251) );
  MUX2X1 U462 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n1195), .Y(n255) );
  MUX2X1 U463 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n1195), .Y(n254) );
  MUX2X1 U464 ( .B(n253), .A(n250), .S(n1175), .Y(n264) );
  MUX2X1 U465 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n1196), .Y(n258) );
  MUX2X1 U466 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n1196), .Y(n257) );
  MUX2X1 U467 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n1196), .Y(n261) );
  MUX2X1 U468 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n1196), .Y(n260) );
  MUX2X1 U469 ( .B(n259), .A(n256), .S(n1175), .Y(n263) );
  MUX2X1 U470 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n1196), .Y(n267) );
  MUX2X1 U471 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n1196), .Y(n266) );
  MUX2X1 U472 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n1196), .Y(n270) );
  MUX2X1 U473 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n1196), .Y(n269) );
  MUX2X1 U474 ( .B(n268), .A(n265), .S(n1175), .Y(n279) );
  MUX2X1 U475 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n1196), .Y(n273) );
  MUX2X1 U476 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n1196), .Y(n272) );
  MUX2X1 U477 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n1196), .Y(n276) );
  MUX2X1 U478 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n1196), .Y(n275) );
  MUX2X1 U479 ( .B(n274), .A(n271), .S(n1175), .Y(n278) );
  MUX2X1 U480 ( .B(n277), .A(n262), .S(n1168), .Y(n643) );
  MUX2X1 U481 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n1197), .Y(n282) );
  MUX2X1 U482 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n1197), .Y(n281) );
  MUX2X1 U483 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n1197), .Y(n285) );
  MUX2X1 U484 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n1197), .Y(n284) );
  MUX2X1 U485 ( .B(n283), .A(n280), .S(n1175), .Y(n294) );
  MUX2X1 U486 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n1197), .Y(n288) );
  MUX2X1 U487 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n1197), .Y(n287) );
  MUX2X1 U488 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n1197), .Y(n291) );
  MUX2X1 U489 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n1197), .Y(n290) );
  MUX2X1 U490 ( .B(n289), .A(n286), .S(n1175), .Y(n293) );
  MUX2X1 U491 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n1197), .Y(n297) );
  MUX2X1 U492 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n1197), .Y(n296) );
  MUX2X1 U493 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n1197), .Y(n300) );
  MUX2X1 U494 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n1197), .Y(n299) );
  MUX2X1 U495 ( .B(n298), .A(n295), .S(n1175), .Y(n309) );
  MUX2X1 U496 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n1194), .Y(n303) );
  MUX2X1 U497 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n1198), .Y(n302) );
  MUX2X1 U498 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n1204), .Y(n306) );
  MUX2X1 U499 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n1198), .Y(n305) );
  MUX2X1 U500 ( .B(n304), .A(n301), .S(n1175), .Y(n308) );
  MUX2X1 U501 ( .B(n307), .A(n292), .S(n1168), .Y(n644) );
  MUX2X1 U502 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n1204), .Y(n312) );
  MUX2X1 U503 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n1194), .Y(n311) );
  MUX2X1 U504 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n1198), .Y(n315) );
  MUX2X1 U505 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n1198), .Y(n314) );
  MUX2X1 U506 ( .B(n313), .A(n310), .S(n1175), .Y(n324) );
  MUX2X1 U507 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n1202), .Y(n318) );
  MUX2X1 U508 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n1201), .Y(n317) );
  MUX2X1 U509 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n1204), .Y(n321) );
  MUX2X1 U510 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n1250), .Y(n320) );
  MUX2X1 U511 ( .B(n319), .A(n316), .S(n1175), .Y(n323) );
  MUX2X1 U512 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n1204), .Y(n327) );
  MUX2X1 U513 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n1194), .Y(n326) );
  MUX2X1 U514 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n1194), .Y(n330) );
  MUX2X1 U515 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n1198), .Y(n329) );
  MUX2X1 U516 ( .B(n328), .A(n325), .S(n1175), .Y(n339) );
  MUX2X1 U517 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n1193), .Y(n333) );
  MUX2X1 U518 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n1195), .Y(n332) );
  MUX2X1 U519 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n1193), .Y(n336) );
  MUX2X1 U520 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n1195), .Y(n335) );
  MUX2X1 U521 ( .B(n334), .A(n331), .S(n1175), .Y(n338) );
  MUX2X1 U522 ( .B(n337), .A(n322), .S(n1168), .Y(n645) );
  MUX2X1 U523 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n1198), .Y(n342) );
  MUX2X1 U524 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n1195), .Y(n341) );
  MUX2X1 U525 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n1204), .Y(n345) );
  MUX2X1 U526 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n1194), .Y(n344) );
  MUX2X1 U527 ( .B(n343), .A(n340), .S(n1174), .Y(n354) );
  MUX2X1 U528 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n1198), .Y(n348) );
  MUX2X1 U529 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n1198), .Y(n347) );
  MUX2X1 U530 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n1198), .Y(n351) );
  MUX2X1 U531 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n1198), .Y(n350) );
  MUX2X1 U532 ( .B(n349), .A(n346), .S(n1174), .Y(n353) );
  MUX2X1 U533 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n1198), .Y(n357) );
  MUX2X1 U534 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n1198), .Y(n356) );
  MUX2X1 U535 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n1198), .Y(n360) );
  MUX2X1 U536 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n1198), .Y(n359) );
  MUX2X1 U537 ( .B(n358), .A(n355), .S(n1174), .Y(n369) );
  MUX2X1 U538 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n1198), .Y(n363) );
  MUX2X1 U539 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n1198), .Y(n362) );
  MUX2X1 U540 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n1198), .Y(n366) );
  MUX2X1 U541 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n1198), .Y(n365) );
  MUX2X1 U542 ( .B(n364), .A(n361), .S(n1174), .Y(n368) );
  MUX2X1 U543 ( .B(n367), .A(n352), .S(n1168), .Y(n646) );
  MUX2X1 U544 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n1204), .Y(n372) );
  MUX2X1 U545 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n1204), .Y(n371) );
  MUX2X1 U546 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n1204), .Y(n375) );
  MUX2X1 U547 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n1194), .Y(n374) );
  MUX2X1 U548 ( .B(n373), .A(n370), .S(n1174), .Y(n384) );
  MUX2X1 U549 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n1194), .Y(n378) );
  MUX2X1 U550 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n1195), .Y(n377) );
  MUX2X1 U551 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n1204), .Y(n381) );
  MUX2X1 U552 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n1194), .Y(n380) );
  MUX2X1 U553 ( .B(n379), .A(n376), .S(n1174), .Y(n383) );
  MUX2X1 U554 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n1194), .Y(n387) );
  MUX2X1 U555 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n1195), .Y(n386) );
  MUX2X1 U556 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n1204), .Y(n390) );
  MUX2X1 U557 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n1195), .Y(n389) );
  MUX2X1 U558 ( .B(n388), .A(n385), .S(n1174), .Y(n399) );
  MUX2X1 U559 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n1199), .Y(n393) );
  MUX2X1 U560 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n1199), .Y(n392) );
  MUX2X1 U561 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n1199), .Y(n396) );
  MUX2X1 U562 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n1199), .Y(n395) );
  MUX2X1 U563 ( .B(n394), .A(n391), .S(n1174), .Y(n398) );
  MUX2X1 U564 ( .B(n397), .A(n382), .S(n1168), .Y(n647) );
  MUX2X1 U565 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n1199), .Y(n402) );
  MUX2X1 U566 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n1199), .Y(n401) );
  MUX2X1 U567 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n1199), .Y(n405) );
  MUX2X1 U568 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n1199), .Y(n404) );
  MUX2X1 U569 ( .B(n403), .A(n400), .S(n1174), .Y(n414) );
  MUX2X1 U570 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n1199), .Y(n408) );
  MUX2X1 U571 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n1199), .Y(n407) );
  MUX2X1 U572 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n1199), .Y(n411) );
  MUX2X1 U573 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n1199), .Y(n410) );
  MUX2X1 U574 ( .B(n409), .A(n406), .S(n1174), .Y(n413) );
  MUX2X1 U575 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n1200), .Y(n417) );
  MUX2X1 U576 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n1200), .Y(n416) );
  MUX2X1 U577 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n1200), .Y(n420) );
  MUX2X1 U578 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n1200), .Y(n419) );
  MUX2X1 U579 ( .B(n418), .A(n415), .S(n1174), .Y(n429) );
  MUX2X1 U580 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n1200), .Y(n423) );
  MUX2X1 U581 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n1200), .Y(n422) );
  MUX2X1 U582 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n1200), .Y(n426) );
  MUX2X1 U583 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n1200), .Y(n425) );
  MUX2X1 U584 ( .B(n424), .A(n421), .S(n1174), .Y(n428) );
  MUX2X1 U585 ( .B(n427), .A(n412), .S(n1168), .Y(n648) );
  MUX2X1 U586 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n1200), .Y(n432) );
  MUX2X1 U587 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n1200), .Y(n431) );
  MUX2X1 U588 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n1200), .Y(n435) );
  MUX2X1 U589 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n1200), .Y(n434) );
  MUX2X1 U590 ( .B(n433), .A(n430), .S(n1173), .Y(n444) );
  MUX2X1 U591 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n1201), .Y(n438) );
  MUX2X1 U592 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n1201), .Y(n437) );
  MUX2X1 U593 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n1201), .Y(n441) );
  MUX2X1 U594 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n1201), .Y(n440) );
  MUX2X1 U595 ( .B(n439), .A(n436), .S(n1173), .Y(n443) );
  MUX2X1 U596 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n1201), .Y(n447) );
  MUX2X1 U597 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n1201), .Y(n446) );
  MUX2X1 U598 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n1201), .Y(n450) );
  MUX2X1 U599 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n1201), .Y(n449) );
  MUX2X1 U600 ( .B(n448), .A(n445), .S(n1173), .Y(n459) );
  MUX2X1 U601 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n1201), .Y(n453) );
  MUX2X1 U602 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n1201), .Y(n452) );
  MUX2X1 U603 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n1201), .Y(n456) );
  MUX2X1 U604 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n1201), .Y(n455) );
  MUX2X1 U605 ( .B(n454), .A(n451), .S(n1173), .Y(n458) );
  MUX2X1 U606 ( .B(n457), .A(n442), .S(n1168), .Y(n649) );
  MUX2X1 U607 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n1202), .Y(n462) );
  MUX2X1 U608 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n1202), .Y(n461) );
  MUX2X1 U609 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n1202), .Y(n465) );
  MUX2X1 U610 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n1202), .Y(n464) );
  MUX2X1 U611 ( .B(n463), .A(n460), .S(n1173), .Y(n474) );
  MUX2X1 U612 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n1202), .Y(n468) );
  MUX2X1 U613 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n1202), .Y(n467) );
  MUX2X1 U614 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n1202), .Y(n471) );
  MUX2X1 U615 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n1202), .Y(n470) );
  MUX2X1 U616 ( .B(n469), .A(n466), .S(n1173), .Y(n473) );
  MUX2X1 U617 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n1202), .Y(n477) );
  MUX2X1 U618 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n1202), .Y(n476) );
  MUX2X1 U619 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n1202), .Y(n480) );
  MUX2X1 U620 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n1202), .Y(n479) );
  MUX2X1 U621 ( .B(n478), .A(n475), .S(n1173), .Y(n489) );
  MUX2X1 U622 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n1203), .Y(n483) );
  MUX2X1 U623 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n1203), .Y(n482) );
  MUX2X1 U624 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n1203), .Y(n486) );
  MUX2X1 U625 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n1203), .Y(n485) );
  MUX2X1 U626 ( .B(n484), .A(n481), .S(n1173), .Y(n488) );
  MUX2X1 U627 ( .B(n487), .A(n472), .S(n1168), .Y(n650) );
  MUX2X1 U628 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n1203), .Y(n492) );
  MUX2X1 U629 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n1203), .Y(n491) );
  MUX2X1 U630 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n1203), .Y(n495) );
  MUX2X1 U631 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n1203), .Y(n494) );
  MUX2X1 U632 ( .B(n493), .A(n490), .S(n1173), .Y(n504) );
  MUX2X1 U633 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n1203), .Y(n498) );
  MUX2X1 U634 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n1203), .Y(n497) );
  MUX2X1 U635 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n1203), .Y(n501) );
  MUX2X1 U636 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n1203), .Y(n500) );
  MUX2X1 U637 ( .B(n499), .A(n496), .S(n1173), .Y(n503) );
  MUX2X1 U638 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n1204), .Y(n507) );
  MUX2X1 U639 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n1204), .Y(n506) );
  MUX2X1 U640 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n1204), .Y(n510) );
  MUX2X1 U641 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n1204), .Y(n509) );
  MUX2X1 U642 ( .B(n508), .A(n505), .S(n1173), .Y(n519) );
  MUX2X1 U643 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n1204), .Y(n513) );
  MUX2X1 U644 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n1204), .Y(n512) );
  MUX2X1 U645 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n1204), .Y(n516) );
  MUX2X1 U646 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n1204), .Y(n515) );
  MUX2X1 U647 ( .B(n514), .A(n511), .S(n1173), .Y(n518) );
  MUX2X1 U648 ( .B(n517), .A(n502), .S(n1168), .Y(n1163) );
  MUX2X1 U649 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n1204), .Y(n522) );
  MUX2X1 U650 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n1204), .Y(n521) );
  MUX2X1 U651 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n1204), .Y(n525) );
  MUX2X1 U652 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n1204), .Y(n524) );
  MUX2X1 U653 ( .B(n523), .A(n520), .S(n1172), .Y(n534) );
  MUX2X1 U654 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n1205), .Y(n528) );
  MUX2X1 U655 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n1205), .Y(n527) );
  MUX2X1 U656 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n1205), .Y(n531) );
  MUX2X1 U657 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n1205), .Y(n530) );
  MUX2X1 U658 ( .B(n529), .A(n526), .S(n1172), .Y(n533) );
  MUX2X1 U659 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n1205), .Y(n537) );
  MUX2X1 U660 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n1205), .Y(n536) );
  MUX2X1 U661 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n1205), .Y(n540) );
  MUX2X1 U662 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n1205), .Y(n539) );
  MUX2X1 U663 ( .B(n538), .A(n535), .S(n1172), .Y(n549) );
  MUX2X1 U664 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n1205), .Y(n543) );
  MUX2X1 U665 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n1205), .Y(n542) );
  MUX2X1 U666 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n1205), .Y(n546) );
  MUX2X1 U667 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n1205), .Y(n545) );
  MUX2X1 U668 ( .B(n544), .A(n541), .S(n1172), .Y(n548) );
  MUX2X1 U669 ( .B(n547), .A(n532), .S(n1168), .Y(n1164) );
  MUX2X1 U670 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n1199), .Y(n552) );
  MUX2X1 U671 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n1194), .Y(n551) );
  MUX2X1 U672 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n1203), .Y(n555) );
  MUX2X1 U673 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n1195), .Y(n554) );
  MUX2X1 U674 ( .B(n553), .A(n550), .S(n1172), .Y(n564) );
  MUX2X1 U675 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n1200), .Y(n558) );
  MUX2X1 U676 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n1204), .Y(n557) );
  MUX2X1 U677 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n1206), .Y(n561) );
  MUX2X1 U678 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n1206), .Y(n560) );
  MUX2X1 U679 ( .B(n559), .A(n556), .S(n1172), .Y(n563) );
  MUX2X1 U680 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n1206), .Y(n567) );
  MUX2X1 U681 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n1206), .Y(n566) );
  MUX2X1 U682 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n1193), .Y(n570) );
  MUX2X1 U683 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n1206), .Y(n569) );
  MUX2X1 U684 ( .B(n568), .A(n565), .S(n1172), .Y(n579) );
  MUX2X1 U685 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n1206), .Y(n573) );
  MUX2X1 U686 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n1206), .Y(n572) );
  MUX2X1 U687 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n1206), .Y(n576) );
  MUX2X1 U688 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n1206), .Y(n575) );
  MUX2X1 U689 ( .B(n574), .A(n571), .S(n1172), .Y(n578) );
  MUX2X1 U690 ( .B(n577), .A(n562), .S(n1168), .Y(n1165) );
  MUX2X1 U691 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n1206), .Y(n582) );
  MUX2X1 U692 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n1206), .Y(n581) );
  MUX2X1 U693 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n1206), .Y(n585) );
  MUX2X1 U694 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n1206), .Y(n584) );
  MUX2X1 U695 ( .B(n583), .A(n580), .S(n1172), .Y(n594) );
  MUX2X1 U696 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n1193), .Y(n588) );
  MUX2X1 U697 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n1202), .Y(n587) );
  MUX2X1 U698 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n1206), .Y(n591) );
  MUX2X1 U699 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n1206), .Y(n590) );
  MUX2X1 U700 ( .B(n589), .A(n586), .S(n1172), .Y(n593) );
  MUX2X1 U701 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n1206), .Y(n597) );
  MUX2X1 U702 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n1206), .Y(n596) );
  MUX2X1 U703 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n1206), .Y(n600) );
  MUX2X1 U704 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n1206), .Y(n599) );
  MUX2X1 U705 ( .B(n598), .A(n595), .S(n1172), .Y(n609) );
  MUX2X1 U706 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n1206), .Y(n603) );
  MUX2X1 U707 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n1206), .Y(n602) );
  MUX2X1 U708 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n1206), .Y(n606) );
  MUX2X1 U709 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n1206), .Y(n605) );
  MUX2X1 U710 ( .B(n604), .A(n601), .S(n1172), .Y(n608) );
  MUX2X1 U711 ( .B(n607), .A(n592), .S(n1168), .Y(n1166) );
  MUX2X1 U712 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n1206), .Y(n612) );
  MUX2X1 U713 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n1206), .Y(n611) );
  MUX2X1 U714 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n1206), .Y(n615) );
  MUX2X1 U715 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n1206), .Y(n614) );
  MUX2X1 U716 ( .B(n613), .A(n610), .S(n1172), .Y(n624) );
  MUX2X1 U717 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n1204), .Y(n618) );
  MUX2X1 U718 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n1200), .Y(n617) );
  MUX2X1 U719 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n1250), .Y(n621) );
  MUX2X1 U720 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n1194), .Y(n620) );
  MUX2X1 U721 ( .B(n619), .A(n616), .S(n1175), .Y(n623) );
  MUX2X1 U722 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n1195), .Y(n627) );
  MUX2X1 U723 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n1196), .Y(n626) );
  MUX2X1 U724 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n1193), .Y(n630) );
  MUX2X1 U725 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n1201), .Y(n629) );
  MUX2X1 U726 ( .B(n628), .A(n625), .S(n1173), .Y(n639) );
  MUX2X1 U727 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n1197), .Y(n633) );
  MUX2X1 U728 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n1195), .Y(n632) );
  MUX2X1 U729 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n1194), .Y(n636) );
  MUX2X1 U730 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n1198), .Y(n635) );
  MUX2X1 U731 ( .B(n634), .A(n631), .S(n1175), .Y(n638) );
  MUX2X1 U732 ( .B(n637), .A(n622), .S(n1168), .Y(n1167) );
  INVX1 U733 ( .A(N12), .Y(n1255) );
  INVX1 U734 ( .A(N11), .Y(n1253) );
  INVX1 U735 ( .A(N10), .Y(n1251) );
  INVX8 U736 ( .A(n1216), .Y(n1211) );
  INVX8 U737 ( .A(n1215), .Y(n1212) );
  INVX8 U738 ( .A(n1215), .Y(n1213) );
  INVX8 U739 ( .A(n36), .Y(n1217) );
  INVX8 U740 ( .A(n36), .Y(n1218) );
  INVX8 U741 ( .A(n37), .Y(n1219) );
  INVX8 U742 ( .A(n37), .Y(n1220) );
  INVX8 U743 ( .A(n38), .Y(n1221) );
  INVX8 U744 ( .A(n38), .Y(n1222) );
  INVX8 U745 ( .A(n39), .Y(n1223) );
  INVX8 U746 ( .A(n39), .Y(n1224) );
  INVX8 U747 ( .A(n40), .Y(n1225) );
  INVX8 U748 ( .A(n40), .Y(n1226) );
  INVX8 U749 ( .A(n41), .Y(n1227) );
  INVX8 U750 ( .A(n41), .Y(n1228) );
  INVX8 U751 ( .A(n42), .Y(n1229) );
  INVX8 U752 ( .A(n42), .Y(n1230) );
  INVX8 U753 ( .A(n43), .Y(n1231) );
  INVX8 U754 ( .A(n43), .Y(n1232) );
  INVX8 U755 ( .A(n44), .Y(n1233) );
  INVX8 U756 ( .A(n44), .Y(n1234) );
  INVX8 U757 ( .A(n45), .Y(n1235) );
  INVX8 U758 ( .A(n45), .Y(n1236) );
  INVX8 U759 ( .A(n46), .Y(n1237) );
  INVX8 U760 ( .A(n46), .Y(n1238) );
  INVX8 U761 ( .A(n61), .Y(n1239) );
  INVX8 U762 ( .A(n61), .Y(n1240) );
  INVX8 U763 ( .A(n62), .Y(n1241) );
  INVX8 U764 ( .A(n62), .Y(n1242) );
  INVX8 U765 ( .A(n63), .Y(n1243) );
  INVX8 U766 ( .A(n63), .Y(n1244) );
  INVX8 U767 ( .A(n64), .Y(n1245) );
  INVX8 U768 ( .A(n64), .Y(n1246) );
  INVX8 U769 ( .A(n65), .Y(n1247) );
  INVX8 U770 ( .A(n65), .Y(n1248) );
  OR2X2 U771 ( .A(write), .B(rst), .Y(n1259) );
  AND2X2 U772 ( .A(n3), .B(N32), .Y(\data_out<0> ) );
  AND2X2 U773 ( .A(n3), .B(N31), .Y(\data_out<1> ) );
  AND2X2 U774 ( .A(n1), .B(N30), .Y(\data_out<2> ) );
  AND2X2 U775 ( .A(n3), .B(N29), .Y(\data_out<3> ) );
  AND2X2 U776 ( .A(n3), .B(N28), .Y(\data_out<4> ) );
  AND2X2 U777 ( .A(n1), .B(N27), .Y(\data_out<5> ) );
  AND2X2 U778 ( .A(n3), .B(N26), .Y(\data_out<6> ) );
  AND2X2 U779 ( .A(n1260), .B(N25), .Y(\data_out<7> ) );
  AND2X2 U780 ( .A(n1), .B(N24), .Y(\data_out<8> ) );
  AND2X2 U781 ( .A(n1), .B(N23), .Y(\data_out<9> ) );
  AND2X2 U782 ( .A(n3), .B(N22), .Y(\data_out<10> ) );
  AND2X2 U783 ( .A(n3), .B(N21), .Y(\data_out<11> ) );
  AND2X2 U784 ( .A(n1260), .B(N20), .Y(\data_out<12> ) );
  AND2X2 U785 ( .A(n1260), .B(N19), .Y(\data_out<13> ) );
  AND2X2 U786 ( .A(n1260), .B(N18), .Y(\data_out<14> ) );
  AND2X2 U787 ( .A(n3), .B(N17), .Y(\data_out<15> ) );
  NAND2X1 U788 ( .A(\mem<31><0> ), .B(n73), .Y(n1261) );
  OAI21X1 U789 ( .A(n72), .B(n1217), .C(n1261), .Y(n2299) );
  NAND2X1 U790 ( .A(\mem<31><1> ), .B(n73), .Y(n1262) );
  OAI21X1 U791 ( .A(n1220), .B(n72), .C(n1262), .Y(n2298) );
  NAND2X1 U792 ( .A(\mem<31><2> ), .B(n73), .Y(n1263) );
  OAI21X1 U793 ( .A(n1222), .B(n72), .C(n1263), .Y(n2297) );
  NAND2X1 U794 ( .A(\mem<31><3> ), .B(n73), .Y(n1264) );
  OAI21X1 U795 ( .A(n1224), .B(n72), .C(n1264), .Y(n2296) );
  NAND2X1 U796 ( .A(\mem<31><4> ), .B(n73), .Y(n1265) );
  OAI21X1 U797 ( .A(n1226), .B(n72), .C(n1265), .Y(n2295) );
  NAND2X1 U798 ( .A(\mem<31><5> ), .B(n73), .Y(n1266) );
  OAI21X1 U799 ( .A(n1228), .B(n72), .C(n1266), .Y(n2294) );
  NAND2X1 U800 ( .A(\mem<31><6> ), .B(n73), .Y(n1267) );
  OAI21X1 U801 ( .A(n1230), .B(n72), .C(n1267), .Y(n2293) );
  NAND2X1 U802 ( .A(\mem<31><7> ), .B(n73), .Y(n1268) );
  OAI21X1 U803 ( .A(n1232), .B(n72), .C(n1268), .Y(n2292) );
  NAND2X1 U804 ( .A(\mem<31><8> ), .B(n73), .Y(n1269) );
  OAI21X1 U805 ( .A(n1234), .B(n72), .C(n1269), .Y(n2291) );
  NAND2X1 U806 ( .A(\mem<31><9> ), .B(n73), .Y(n1270) );
  OAI21X1 U807 ( .A(n1236), .B(n72), .C(n1270), .Y(n2290) );
  NAND2X1 U808 ( .A(\mem<31><10> ), .B(n73), .Y(n1271) );
  OAI21X1 U809 ( .A(n1238), .B(n72), .C(n1271), .Y(n2289) );
  NAND2X1 U810 ( .A(\mem<31><11> ), .B(n73), .Y(n1272) );
  OAI21X1 U811 ( .A(n1240), .B(n72), .C(n1272), .Y(n2288) );
  NAND2X1 U812 ( .A(\mem<31><12> ), .B(n73), .Y(n1273) );
  OAI21X1 U813 ( .A(n1242), .B(n72), .C(n1273), .Y(n2287) );
  NAND2X1 U814 ( .A(\mem<31><13> ), .B(n73), .Y(n1274) );
  OAI21X1 U815 ( .A(n1244), .B(n72), .C(n1274), .Y(n2286) );
  NAND2X1 U816 ( .A(\mem<31><14> ), .B(n73), .Y(n1275) );
  OAI21X1 U817 ( .A(n1246), .B(n72), .C(n1275), .Y(n2285) );
  NAND2X1 U818 ( .A(\mem<31><15> ), .B(n73), .Y(n1276) );
  OAI21X1 U819 ( .A(n1248), .B(n72), .C(n1276), .Y(n2284) );
  NAND2X1 U820 ( .A(\mem<30><0> ), .B(n76), .Y(n1277) );
  OAI21X1 U821 ( .A(n75), .B(n1217), .C(n1277), .Y(n2283) );
  NAND2X1 U822 ( .A(\mem<30><1> ), .B(n76), .Y(n1278) );
  OAI21X1 U823 ( .A(n75), .B(n1220), .C(n1278), .Y(n2282) );
  NAND2X1 U824 ( .A(\mem<30><2> ), .B(n76), .Y(n1279) );
  OAI21X1 U825 ( .A(n75), .B(n1222), .C(n1279), .Y(n2281) );
  NAND2X1 U826 ( .A(\mem<30><3> ), .B(n76), .Y(n1280) );
  OAI21X1 U827 ( .A(n75), .B(n1224), .C(n1280), .Y(n2280) );
  NAND2X1 U828 ( .A(\mem<30><4> ), .B(n76), .Y(n1281) );
  OAI21X1 U829 ( .A(n75), .B(n1226), .C(n1281), .Y(n2279) );
  NAND2X1 U830 ( .A(\mem<30><5> ), .B(n76), .Y(n1282) );
  OAI21X1 U831 ( .A(n75), .B(n1228), .C(n1282), .Y(n2278) );
  NAND2X1 U832 ( .A(\mem<30><6> ), .B(n76), .Y(n1283) );
  OAI21X1 U833 ( .A(n75), .B(n1230), .C(n1283), .Y(n2277) );
  NAND2X1 U834 ( .A(\mem<30><7> ), .B(n76), .Y(n1284) );
  OAI21X1 U835 ( .A(n75), .B(n1232), .C(n1284), .Y(n2276) );
  NAND2X1 U836 ( .A(\mem<30><8> ), .B(n76), .Y(n1285) );
  OAI21X1 U837 ( .A(n75), .B(n1233), .C(n1285), .Y(n2275) );
  NAND2X1 U838 ( .A(\mem<30><9> ), .B(n76), .Y(n1286) );
  OAI21X1 U839 ( .A(n75), .B(n1235), .C(n1286), .Y(n2274) );
  NAND2X1 U840 ( .A(\mem<30><10> ), .B(n76), .Y(n1287) );
  OAI21X1 U841 ( .A(n75), .B(n1237), .C(n1287), .Y(n2273) );
  NAND2X1 U842 ( .A(\mem<30><11> ), .B(n76), .Y(n1288) );
  OAI21X1 U843 ( .A(n75), .B(n1239), .C(n1288), .Y(n2272) );
  NAND2X1 U844 ( .A(\mem<30><12> ), .B(n76), .Y(n1289) );
  OAI21X1 U845 ( .A(n75), .B(n1241), .C(n1289), .Y(n2271) );
  NAND2X1 U846 ( .A(\mem<30><13> ), .B(n76), .Y(n1290) );
  OAI21X1 U847 ( .A(n75), .B(n1243), .C(n1290), .Y(n2270) );
  NAND2X1 U848 ( .A(\mem<30><14> ), .B(n76), .Y(n1291) );
  OAI21X1 U849 ( .A(n75), .B(n1245), .C(n1291), .Y(n2269) );
  NAND2X1 U850 ( .A(\mem<30><15> ), .B(n76), .Y(n1292) );
  OAI21X1 U851 ( .A(n75), .B(n1247), .C(n1292), .Y(n2268) );
  NAND3X1 U852 ( .A(n1250), .B(n1254), .C(n1253), .Y(n1293) );
  NAND2X1 U853 ( .A(\mem<29><0> ), .B(n79), .Y(n1294) );
  OAI21X1 U854 ( .A(n78), .B(n1217), .C(n1294), .Y(n2267) );
  NAND2X1 U855 ( .A(\mem<29><1> ), .B(n79), .Y(n1295) );
  OAI21X1 U856 ( .A(n78), .B(n1219), .C(n1295), .Y(n2266) );
  NAND2X1 U857 ( .A(\mem<29><2> ), .B(n79), .Y(n1296) );
  OAI21X1 U858 ( .A(n78), .B(n1221), .C(n1296), .Y(n2265) );
  NAND2X1 U859 ( .A(\mem<29><3> ), .B(n79), .Y(n1297) );
  OAI21X1 U860 ( .A(n78), .B(n1223), .C(n1297), .Y(n2264) );
  NAND2X1 U861 ( .A(\mem<29><4> ), .B(n79), .Y(n1298) );
  OAI21X1 U862 ( .A(n78), .B(n1225), .C(n1298), .Y(n2263) );
  NAND2X1 U863 ( .A(\mem<29><5> ), .B(n79), .Y(n1299) );
  OAI21X1 U864 ( .A(n78), .B(n1227), .C(n1299), .Y(n2262) );
  NAND2X1 U865 ( .A(\mem<29><6> ), .B(n79), .Y(n1300) );
  OAI21X1 U866 ( .A(n78), .B(n1229), .C(n1300), .Y(n2261) );
  NAND2X1 U867 ( .A(\mem<29><7> ), .B(n79), .Y(n1301) );
  OAI21X1 U868 ( .A(n78), .B(n1231), .C(n1301), .Y(n2260) );
  NAND2X1 U869 ( .A(\mem<29><8> ), .B(n79), .Y(n1302) );
  OAI21X1 U870 ( .A(n78), .B(n1234), .C(n1302), .Y(n2259) );
  NAND2X1 U871 ( .A(\mem<29><9> ), .B(n79), .Y(n1303) );
  OAI21X1 U872 ( .A(n78), .B(n1236), .C(n1303), .Y(n2258) );
  NAND2X1 U873 ( .A(\mem<29><10> ), .B(n79), .Y(n1304) );
  OAI21X1 U874 ( .A(n78), .B(n1238), .C(n1304), .Y(n2257) );
  NAND2X1 U875 ( .A(\mem<29><11> ), .B(n79), .Y(n1305) );
  OAI21X1 U876 ( .A(n78), .B(n1240), .C(n1305), .Y(n2256) );
  NAND2X1 U877 ( .A(\mem<29><12> ), .B(n79), .Y(n1306) );
  OAI21X1 U878 ( .A(n78), .B(n1242), .C(n1306), .Y(n2255) );
  NAND2X1 U879 ( .A(\mem<29><13> ), .B(n79), .Y(n1307) );
  OAI21X1 U880 ( .A(n78), .B(n1244), .C(n1307), .Y(n2254) );
  NAND2X1 U881 ( .A(\mem<29><14> ), .B(n79), .Y(n1308) );
  OAI21X1 U882 ( .A(n78), .B(n1246), .C(n1308), .Y(n2253) );
  NAND2X1 U883 ( .A(\mem<29><15> ), .B(n79), .Y(n1309) );
  OAI21X1 U884 ( .A(n78), .B(n1248), .C(n1309), .Y(n2252) );
  NAND3X1 U885 ( .A(n1254), .B(n1253), .C(n1251), .Y(n1310) );
  NAND2X1 U886 ( .A(\mem<28><0> ), .B(n82), .Y(n1311) );
  OAI21X1 U887 ( .A(n81), .B(n1217), .C(n1311), .Y(n2251) );
  NAND2X1 U888 ( .A(\mem<28><1> ), .B(n82), .Y(n1312) );
  OAI21X1 U889 ( .A(n81), .B(n1220), .C(n1312), .Y(n2250) );
  NAND2X1 U890 ( .A(\mem<28><2> ), .B(n82), .Y(n1313) );
  OAI21X1 U891 ( .A(n81), .B(n1222), .C(n1313), .Y(n2249) );
  NAND2X1 U892 ( .A(\mem<28><3> ), .B(n82), .Y(n1314) );
  OAI21X1 U893 ( .A(n81), .B(n1224), .C(n1314), .Y(n2248) );
  NAND2X1 U894 ( .A(\mem<28><4> ), .B(n82), .Y(n1315) );
  OAI21X1 U895 ( .A(n81), .B(n1226), .C(n1315), .Y(n2247) );
  NAND2X1 U896 ( .A(\mem<28><5> ), .B(n82), .Y(n1316) );
  OAI21X1 U897 ( .A(n81), .B(n1228), .C(n1316), .Y(n2246) );
  NAND2X1 U898 ( .A(\mem<28><6> ), .B(n82), .Y(n1317) );
  OAI21X1 U899 ( .A(n81), .B(n1230), .C(n1317), .Y(n2245) );
  NAND2X1 U900 ( .A(\mem<28><7> ), .B(n82), .Y(n1318) );
  OAI21X1 U901 ( .A(n81), .B(n1232), .C(n1318), .Y(n2244) );
  NAND2X1 U902 ( .A(\mem<28><8> ), .B(n82), .Y(n1319) );
  OAI21X1 U903 ( .A(n81), .B(n1233), .C(n1319), .Y(n2243) );
  NAND2X1 U904 ( .A(\mem<28><9> ), .B(n82), .Y(n1320) );
  OAI21X1 U905 ( .A(n81), .B(n1235), .C(n1320), .Y(n2242) );
  NAND2X1 U906 ( .A(\mem<28><10> ), .B(n82), .Y(n1321) );
  OAI21X1 U907 ( .A(n81), .B(n1237), .C(n1321), .Y(n2241) );
  NAND2X1 U908 ( .A(\mem<28><11> ), .B(n82), .Y(n1322) );
  OAI21X1 U909 ( .A(n81), .B(n1239), .C(n1322), .Y(n2240) );
  NAND2X1 U910 ( .A(\mem<28><12> ), .B(n82), .Y(n1323) );
  OAI21X1 U911 ( .A(n81), .B(n1241), .C(n1323), .Y(n2239) );
  NAND2X1 U912 ( .A(\mem<28><13> ), .B(n82), .Y(n1324) );
  OAI21X1 U913 ( .A(n81), .B(n1243), .C(n1324), .Y(n2238) );
  NAND2X1 U914 ( .A(\mem<28><14> ), .B(n82), .Y(n1325) );
  OAI21X1 U915 ( .A(n81), .B(n1245), .C(n1325), .Y(n2237) );
  NAND2X1 U916 ( .A(\mem<28><15> ), .B(n82), .Y(n1326) );
  OAI21X1 U917 ( .A(n81), .B(n1247), .C(n1326), .Y(n2236) );
  NAND3X1 U918 ( .A(n1250), .B(n1252), .C(n1255), .Y(n1327) );
  NAND2X1 U919 ( .A(\mem<27><0> ), .B(n85), .Y(n1328) );
  OAI21X1 U920 ( .A(n84), .B(n1217), .C(n1328), .Y(n2235) );
  NAND2X1 U921 ( .A(\mem<27><1> ), .B(n85), .Y(n1329) );
  OAI21X1 U922 ( .A(n84), .B(n1219), .C(n1329), .Y(n2234) );
  NAND2X1 U923 ( .A(\mem<27><2> ), .B(n85), .Y(n1330) );
  OAI21X1 U924 ( .A(n84), .B(n1221), .C(n1330), .Y(n2233) );
  NAND2X1 U925 ( .A(\mem<27><3> ), .B(n85), .Y(n1331) );
  OAI21X1 U926 ( .A(n84), .B(n1223), .C(n1331), .Y(n2232) );
  NAND2X1 U927 ( .A(\mem<27><4> ), .B(n85), .Y(n1332) );
  OAI21X1 U928 ( .A(n84), .B(n1225), .C(n1332), .Y(n2231) );
  NAND2X1 U929 ( .A(\mem<27><5> ), .B(n85), .Y(n1333) );
  OAI21X1 U930 ( .A(n84), .B(n1227), .C(n1333), .Y(n2230) );
  NAND2X1 U931 ( .A(\mem<27><6> ), .B(n85), .Y(n1334) );
  OAI21X1 U932 ( .A(n84), .B(n1229), .C(n1334), .Y(n2229) );
  NAND2X1 U933 ( .A(\mem<27><7> ), .B(n85), .Y(n1335) );
  OAI21X1 U934 ( .A(n84), .B(n1231), .C(n1335), .Y(n2228) );
  NAND2X1 U935 ( .A(\mem<27><8> ), .B(n85), .Y(n1336) );
  OAI21X1 U936 ( .A(n84), .B(n1234), .C(n1336), .Y(n2227) );
  NAND2X1 U937 ( .A(\mem<27><9> ), .B(n85), .Y(n1337) );
  OAI21X1 U938 ( .A(n84), .B(n1236), .C(n1337), .Y(n2226) );
  NAND2X1 U939 ( .A(\mem<27><10> ), .B(n85), .Y(n1338) );
  OAI21X1 U940 ( .A(n84), .B(n1238), .C(n1338), .Y(n2225) );
  NAND2X1 U941 ( .A(\mem<27><11> ), .B(n85), .Y(n1339) );
  OAI21X1 U942 ( .A(n84), .B(n1240), .C(n1339), .Y(n2224) );
  NAND2X1 U943 ( .A(\mem<27><12> ), .B(n85), .Y(n1340) );
  OAI21X1 U944 ( .A(n84), .B(n1242), .C(n1340), .Y(n2223) );
  NAND2X1 U945 ( .A(\mem<27><13> ), .B(n85), .Y(n1341) );
  OAI21X1 U946 ( .A(n84), .B(n1244), .C(n1341), .Y(n2222) );
  NAND2X1 U947 ( .A(\mem<27><14> ), .B(n85), .Y(n1342) );
  OAI21X1 U948 ( .A(n84), .B(n1246), .C(n1342), .Y(n2221) );
  NAND2X1 U949 ( .A(\mem<27><15> ), .B(n85), .Y(n1343) );
  OAI21X1 U950 ( .A(n84), .B(n1248), .C(n1343), .Y(n2220) );
  NAND3X1 U951 ( .A(n1255), .B(n1252), .C(n1251), .Y(n1344) );
  NAND2X1 U952 ( .A(\mem<26><0> ), .B(n88), .Y(n1345) );
  OAI21X1 U953 ( .A(n87), .B(n1217), .C(n1345), .Y(n2219) );
  NAND2X1 U954 ( .A(\mem<26><1> ), .B(n88), .Y(n1346) );
  OAI21X1 U955 ( .A(n87), .B(n1220), .C(n1346), .Y(n2218) );
  NAND2X1 U956 ( .A(\mem<26><2> ), .B(n88), .Y(n1347) );
  OAI21X1 U957 ( .A(n87), .B(n1222), .C(n1347), .Y(n2217) );
  NAND2X1 U958 ( .A(\mem<26><3> ), .B(n88), .Y(n1348) );
  OAI21X1 U959 ( .A(n87), .B(n1224), .C(n1348), .Y(n2216) );
  NAND2X1 U960 ( .A(\mem<26><4> ), .B(n88), .Y(n1349) );
  OAI21X1 U961 ( .A(n87), .B(n1226), .C(n1349), .Y(n2215) );
  NAND2X1 U962 ( .A(\mem<26><5> ), .B(n88), .Y(n1350) );
  OAI21X1 U963 ( .A(n87), .B(n1228), .C(n1350), .Y(n2214) );
  NAND2X1 U964 ( .A(\mem<26><6> ), .B(n88), .Y(n1351) );
  OAI21X1 U965 ( .A(n87), .B(n1230), .C(n1351), .Y(n2213) );
  NAND2X1 U966 ( .A(\mem<26><7> ), .B(n88), .Y(n1352) );
  OAI21X1 U967 ( .A(n87), .B(n1232), .C(n1352), .Y(n2212) );
  NAND2X1 U968 ( .A(\mem<26><8> ), .B(n88), .Y(n1353) );
  OAI21X1 U969 ( .A(n87), .B(n1233), .C(n1353), .Y(n2211) );
  NAND2X1 U970 ( .A(\mem<26><9> ), .B(n88), .Y(n1354) );
  OAI21X1 U971 ( .A(n87), .B(n1235), .C(n1354), .Y(n2210) );
  NAND2X1 U972 ( .A(\mem<26><10> ), .B(n88), .Y(n1355) );
  OAI21X1 U973 ( .A(n87), .B(n1237), .C(n1355), .Y(n2209) );
  NAND2X1 U974 ( .A(\mem<26><11> ), .B(n88), .Y(n1356) );
  OAI21X1 U975 ( .A(n87), .B(n1239), .C(n1356), .Y(n2208) );
  NAND2X1 U976 ( .A(\mem<26><12> ), .B(n88), .Y(n1357) );
  OAI21X1 U977 ( .A(n87), .B(n1241), .C(n1357), .Y(n2207) );
  NAND2X1 U978 ( .A(\mem<26><13> ), .B(n88), .Y(n1358) );
  OAI21X1 U979 ( .A(n87), .B(n1243), .C(n1358), .Y(n2206) );
  NAND2X1 U980 ( .A(\mem<26><14> ), .B(n88), .Y(n1359) );
  OAI21X1 U981 ( .A(n87), .B(n1245), .C(n1359), .Y(n2205) );
  NAND2X1 U982 ( .A(\mem<26><15> ), .B(n88), .Y(n1360) );
  OAI21X1 U983 ( .A(n87), .B(n1247), .C(n1360), .Y(n2204) );
  NAND3X1 U984 ( .A(n1250), .B(n1255), .C(n1253), .Y(n1361) );
  NAND2X1 U985 ( .A(\mem<25><0> ), .B(n91), .Y(n1362) );
  OAI21X1 U986 ( .A(n90), .B(n1217), .C(n1362), .Y(n2203) );
  NAND2X1 U987 ( .A(\mem<25><1> ), .B(n91), .Y(n1363) );
  OAI21X1 U988 ( .A(n90), .B(n1219), .C(n1363), .Y(n2202) );
  NAND2X1 U989 ( .A(\mem<25><2> ), .B(n91), .Y(n1364) );
  OAI21X1 U990 ( .A(n90), .B(n1221), .C(n1364), .Y(n2201) );
  NAND2X1 U991 ( .A(\mem<25><3> ), .B(n91), .Y(n1365) );
  OAI21X1 U992 ( .A(n90), .B(n1223), .C(n1365), .Y(n2200) );
  NAND2X1 U993 ( .A(\mem<25><4> ), .B(n91), .Y(n1366) );
  OAI21X1 U994 ( .A(n90), .B(n1225), .C(n1366), .Y(n2199) );
  NAND2X1 U995 ( .A(\mem<25><5> ), .B(n91), .Y(n1367) );
  OAI21X1 U996 ( .A(n90), .B(n1227), .C(n1367), .Y(n2198) );
  NAND2X1 U997 ( .A(\mem<25><6> ), .B(n91), .Y(n1368) );
  OAI21X1 U998 ( .A(n90), .B(n1229), .C(n1368), .Y(n2197) );
  NAND2X1 U999 ( .A(\mem<25><7> ), .B(n91), .Y(n1369) );
  OAI21X1 U1000 ( .A(n90), .B(n1231), .C(n1369), .Y(n2196) );
  NAND2X1 U1001 ( .A(\mem<25><8> ), .B(n91), .Y(n1370) );
  OAI21X1 U1002 ( .A(n90), .B(n1234), .C(n1370), .Y(n2195) );
  NAND2X1 U1003 ( .A(\mem<25><9> ), .B(n91), .Y(n1371) );
  OAI21X1 U1004 ( .A(n90), .B(n1236), .C(n1371), .Y(n2194) );
  NAND2X1 U1005 ( .A(\mem<25><10> ), .B(n91), .Y(n1372) );
  OAI21X1 U1006 ( .A(n90), .B(n1238), .C(n1372), .Y(n2193) );
  NAND2X1 U1007 ( .A(\mem<25><11> ), .B(n91), .Y(n1373) );
  OAI21X1 U1008 ( .A(n90), .B(n1240), .C(n1373), .Y(n2192) );
  NAND2X1 U1009 ( .A(\mem<25><12> ), .B(n91), .Y(n1374) );
  OAI21X1 U1010 ( .A(n90), .B(n1242), .C(n1374), .Y(n2191) );
  NAND2X1 U1011 ( .A(\mem<25><13> ), .B(n91), .Y(n1375) );
  OAI21X1 U1012 ( .A(n90), .B(n1244), .C(n1375), .Y(n2190) );
  NAND2X1 U1013 ( .A(\mem<25><14> ), .B(n91), .Y(n1376) );
  OAI21X1 U1014 ( .A(n90), .B(n1246), .C(n1376), .Y(n2189) );
  NAND2X1 U1015 ( .A(\mem<25><15> ), .B(n91), .Y(n1377) );
  OAI21X1 U1016 ( .A(n90), .B(n1248), .C(n1377), .Y(n2188) );
  NOR3X1 U1017 ( .A(n1250), .B(n1252), .C(n1254), .Y(n1771) );
  NAND2X1 U1018 ( .A(\mem<24><0> ), .B(n92), .Y(n1378) );
  OAI21X1 U1019 ( .A(n1208), .B(n1217), .C(n1378), .Y(n2187) );
  NAND2X1 U1020 ( .A(\mem<24><1> ), .B(n92), .Y(n1379) );
  OAI21X1 U1021 ( .A(n1208), .B(n1219), .C(n1379), .Y(n2186) );
  NAND2X1 U1022 ( .A(\mem<24><2> ), .B(n92), .Y(n1380) );
  OAI21X1 U1023 ( .A(n1208), .B(n1221), .C(n1380), .Y(n2185) );
  NAND2X1 U1024 ( .A(\mem<24><3> ), .B(n92), .Y(n1381) );
  OAI21X1 U1025 ( .A(n1208), .B(n1223), .C(n1381), .Y(n2184) );
  NAND2X1 U1026 ( .A(\mem<24><4> ), .B(n92), .Y(n1382) );
  OAI21X1 U1027 ( .A(n1208), .B(n1225), .C(n1382), .Y(n2183) );
  NAND2X1 U1028 ( .A(\mem<24><5> ), .B(n92), .Y(n1383) );
  OAI21X1 U1029 ( .A(n1208), .B(n1227), .C(n1383), .Y(n2182) );
  NAND2X1 U1030 ( .A(\mem<24><6> ), .B(n92), .Y(n1384) );
  OAI21X1 U1031 ( .A(n1208), .B(n1229), .C(n1384), .Y(n2181) );
  NAND2X1 U1032 ( .A(\mem<24><7> ), .B(n92), .Y(n1385) );
  OAI21X1 U1033 ( .A(n1208), .B(n1231), .C(n1385), .Y(n2180) );
  NAND2X1 U1034 ( .A(\mem<24><8> ), .B(n92), .Y(n1386) );
  OAI21X1 U1035 ( .A(n1208), .B(n1233), .C(n1386), .Y(n2179) );
  NAND2X1 U1036 ( .A(\mem<24><9> ), .B(n92), .Y(n1387) );
  OAI21X1 U1037 ( .A(n1208), .B(n1235), .C(n1387), .Y(n2178) );
  NAND2X1 U1038 ( .A(\mem<24><10> ), .B(n92), .Y(n1388) );
  OAI21X1 U1039 ( .A(n1208), .B(n1237), .C(n1388), .Y(n2177) );
  NAND2X1 U1040 ( .A(\mem<24><11> ), .B(n92), .Y(n1389) );
  OAI21X1 U1041 ( .A(n1208), .B(n1239), .C(n1389), .Y(n2176) );
  NAND2X1 U1042 ( .A(\mem<24><12> ), .B(n92), .Y(n1390) );
  OAI21X1 U1043 ( .A(n1208), .B(n1241), .C(n1390), .Y(n2175) );
  NAND2X1 U1044 ( .A(\mem<24><13> ), .B(n92), .Y(n1391) );
  OAI21X1 U1045 ( .A(n1208), .B(n1243), .C(n1391), .Y(n2174) );
  NAND2X1 U1046 ( .A(\mem<24><14> ), .B(n92), .Y(n1392) );
  OAI21X1 U1047 ( .A(n1208), .B(n1245), .C(n1392), .Y(n2173) );
  NAND2X1 U1048 ( .A(\mem<24><15> ), .B(n92), .Y(n1393) );
  OAI21X1 U1049 ( .A(n1208), .B(n1247), .C(n1393), .Y(n2172) );
  NAND2X1 U1050 ( .A(\mem<23><0> ), .B(n95), .Y(n1394) );
  OAI21X1 U1051 ( .A(n94), .B(n1217), .C(n1394), .Y(n2171) );
  NAND2X1 U1052 ( .A(\mem<23><1> ), .B(n95), .Y(n1395) );
  OAI21X1 U1053 ( .A(n94), .B(n1220), .C(n1395), .Y(n2170) );
  NAND2X1 U1054 ( .A(\mem<23><2> ), .B(n95), .Y(n1396) );
  OAI21X1 U1055 ( .A(n94), .B(n1222), .C(n1396), .Y(n2169) );
  NAND2X1 U1056 ( .A(\mem<23><3> ), .B(n95), .Y(n1397) );
  OAI21X1 U1057 ( .A(n94), .B(n1224), .C(n1397), .Y(n2168) );
  NAND2X1 U1058 ( .A(\mem<23><4> ), .B(n95), .Y(n1398) );
  OAI21X1 U1059 ( .A(n94), .B(n1226), .C(n1398), .Y(n2167) );
  NAND2X1 U1060 ( .A(\mem<23><5> ), .B(n95), .Y(n1399) );
  OAI21X1 U1061 ( .A(n94), .B(n1228), .C(n1399), .Y(n2166) );
  NAND2X1 U1062 ( .A(\mem<23><6> ), .B(n95), .Y(n1400) );
  OAI21X1 U1063 ( .A(n94), .B(n1230), .C(n1400), .Y(n2165) );
  NAND2X1 U1064 ( .A(\mem<23><7> ), .B(n95), .Y(n1401) );
  OAI21X1 U1065 ( .A(n94), .B(n1232), .C(n1401), .Y(n2164) );
  NAND2X1 U1066 ( .A(\mem<23><8> ), .B(n95), .Y(n1402) );
  OAI21X1 U1067 ( .A(n94), .B(n1234), .C(n1402), .Y(n2163) );
  NAND2X1 U1068 ( .A(\mem<23><9> ), .B(n95), .Y(n1403) );
  OAI21X1 U1069 ( .A(n94), .B(n1236), .C(n1403), .Y(n2162) );
  NAND2X1 U1070 ( .A(\mem<23><10> ), .B(n95), .Y(n1404) );
  OAI21X1 U1071 ( .A(n94), .B(n1238), .C(n1404), .Y(n2161) );
  NAND2X1 U1072 ( .A(\mem<23><11> ), .B(n95), .Y(n1405) );
  OAI21X1 U1073 ( .A(n94), .B(n1240), .C(n1405), .Y(n2160) );
  NAND2X1 U1074 ( .A(\mem<23><12> ), .B(n95), .Y(n1406) );
  OAI21X1 U1075 ( .A(n94), .B(n1242), .C(n1406), .Y(n2159) );
  NAND2X1 U1076 ( .A(\mem<23><13> ), .B(n95), .Y(n1407) );
  OAI21X1 U1077 ( .A(n94), .B(n1244), .C(n1407), .Y(n2158) );
  NAND2X1 U1078 ( .A(\mem<23><14> ), .B(n95), .Y(n1408) );
  OAI21X1 U1079 ( .A(n94), .B(n1246), .C(n1408), .Y(n2157) );
  NAND2X1 U1080 ( .A(\mem<23><15> ), .B(n95), .Y(n1409) );
  OAI21X1 U1081 ( .A(n94), .B(n1248), .C(n1409), .Y(n2156) );
  NAND2X1 U1082 ( .A(\mem<22><0> ), .B(n98), .Y(n1410) );
  OAI21X1 U1083 ( .A(n97), .B(n1217), .C(n1410), .Y(n2155) );
  NAND2X1 U1084 ( .A(\mem<22><1> ), .B(n98), .Y(n1411) );
  OAI21X1 U1085 ( .A(n97), .B(n1220), .C(n1411), .Y(n2154) );
  NAND2X1 U1086 ( .A(\mem<22><2> ), .B(n98), .Y(n1412) );
  OAI21X1 U1087 ( .A(n97), .B(n1222), .C(n1412), .Y(n2153) );
  NAND2X1 U1088 ( .A(\mem<22><3> ), .B(n98), .Y(n1413) );
  OAI21X1 U1089 ( .A(n97), .B(n1224), .C(n1413), .Y(n2152) );
  NAND2X1 U1090 ( .A(\mem<22><4> ), .B(n98), .Y(n1414) );
  OAI21X1 U1091 ( .A(n97), .B(n1226), .C(n1414), .Y(n2151) );
  NAND2X1 U1092 ( .A(\mem<22><5> ), .B(n98), .Y(n1415) );
  OAI21X1 U1093 ( .A(n97), .B(n1228), .C(n1415), .Y(n2150) );
  NAND2X1 U1094 ( .A(\mem<22><6> ), .B(n98), .Y(n1416) );
  OAI21X1 U1095 ( .A(n97), .B(n1230), .C(n1416), .Y(n2149) );
  NAND2X1 U1096 ( .A(\mem<22><7> ), .B(n98), .Y(n1417) );
  OAI21X1 U1097 ( .A(n97), .B(n1232), .C(n1417), .Y(n2148) );
  NAND2X1 U1098 ( .A(\mem<22><8> ), .B(n98), .Y(n1418) );
  OAI21X1 U1099 ( .A(n97), .B(n1234), .C(n1418), .Y(n2147) );
  NAND2X1 U1100 ( .A(\mem<22><9> ), .B(n98), .Y(n1419) );
  OAI21X1 U1101 ( .A(n97), .B(n1236), .C(n1419), .Y(n2146) );
  NAND2X1 U1102 ( .A(\mem<22><10> ), .B(n98), .Y(n1420) );
  OAI21X1 U1103 ( .A(n97), .B(n1238), .C(n1420), .Y(n2145) );
  NAND2X1 U1104 ( .A(\mem<22><11> ), .B(n98), .Y(n1421) );
  OAI21X1 U1105 ( .A(n97), .B(n1240), .C(n1421), .Y(n2144) );
  NAND2X1 U1106 ( .A(\mem<22><12> ), .B(n98), .Y(n1422) );
  OAI21X1 U1107 ( .A(n97), .B(n1242), .C(n1422), .Y(n2143) );
  NAND2X1 U1108 ( .A(\mem<22><13> ), .B(n98), .Y(n1423) );
  OAI21X1 U1109 ( .A(n97), .B(n1244), .C(n1423), .Y(n2142) );
  NAND2X1 U1110 ( .A(\mem<22><14> ), .B(n98), .Y(n1424) );
  OAI21X1 U1111 ( .A(n97), .B(n1246), .C(n1424), .Y(n2141) );
  NAND2X1 U1112 ( .A(\mem<22><15> ), .B(n98), .Y(n1425) );
  OAI21X1 U1113 ( .A(n97), .B(n1248), .C(n1425), .Y(n2140) );
  NAND2X1 U1114 ( .A(\mem<21><0> ), .B(n101), .Y(n1426) );
  OAI21X1 U1115 ( .A(n100), .B(n1217), .C(n1426), .Y(n2139) );
  NAND2X1 U1116 ( .A(\mem<21><1> ), .B(n101), .Y(n1427) );
  OAI21X1 U1117 ( .A(n100), .B(n1220), .C(n1427), .Y(n2138) );
  NAND2X1 U1118 ( .A(\mem<21><2> ), .B(n101), .Y(n1428) );
  OAI21X1 U1119 ( .A(n100), .B(n1222), .C(n1428), .Y(n2137) );
  NAND2X1 U1120 ( .A(\mem<21><3> ), .B(n101), .Y(n1429) );
  OAI21X1 U1121 ( .A(n100), .B(n1224), .C(n1429), .Y(n2136) );
  NAND2X1 U1122 ( .A(\mem<21><4> ), .B(n101), .Y(n1430) );
  OAI21X1 U1123 ( .A(n100), .B(n1226), .C(n1430), .Y(n2135) );
  NAND2X1 U1124 ( .A(\mem<21><5> ), .B(n101), .Y(n1431) );
  OAI21X1 U1125 ( .A(n100), .B(n1228), .C(n1431), .Y(n2134) );
  NAND2X1 U1126 ( .A(\mem<21><6> ), .B(n101), .Y(n1432) );
  OAI21X1 U1127 ( .A(n100), .B(n1230), .C(n1432), .Y(n2133) );
  NAND2X1 U1128 ( .A(\mem<21><7> ), .B(n101), .Y(n1433) );
  OAI21X1 U1129 ( .A(n100), .B(n1232), .C(n1433), .Y(n2132) );
  NAND2X1 U1130 ( .A(\mem<21><8> ), .B(n101), .Y(n1434) );
  OAI21X1 U1131 ( .A(n100), .B(n1234), .C(n1434), .Y(n2131) );
  NAND2X1 U1132 ( .A(\mem<21><9> ), .B(n101), .Y(n1435) );
  OAI21X1 U1133 ( .A(n100), .B(n1236), .C(n1435), .Y(n2130) );
  NAND2X1 U1134 ( .A(\mem<21><10> ), .B(n101), .Y(n1436) );
  OAI21X1 U1135 ( .A(n100), .B(n1238), .C(n1436), .Y(n2129) );
  NAND2X1 U1136 ( .A(\mem<21><11> ), .B(n101), .Y(n1437) );
  OAI21X1 U1137 ( .A(n100), .B(n1240), .C(n1437), .Y(n2128) );
  NAND2X1 U1138 ( .A(\mem<21><12> ), .B(n101), .Y(n1438) );
  OAI21X1 U1139 ( .A(n100), .B(n1242), .C(n1438), .Y(n2127) );
  NAND2X1 U1140 ( .A(\mem<21><13> ), .B(n101), .Y(n1439) );
  OAI21X1 U1141 ( .A(n100), .B(n1244), .C(n1439), .Y(n2126) );
  NAND2X1 U1142 ( .A(\mem<21><14> ), .B(n101), .Y(n1440) );
  OAI21X1 U1143 ( .A(n100), .B(n1246), .C(n1440), .Y(n2125) );
  NAND2X1 U1144 ( .A(\mem<21><15> ), .B(n101), .Y(n1441) );
  OAI21X1 U1145 ( .A(n100), .B(n1248), .C(n1441), .Y(n2124) );
  NAND2X1 U1146 ( .A(\mem<20><0> ), .B(n104), .Y(n1442) );
  OAI21X1 U1147 ( .A(n103), .B(n1217), .C(n1442), .Y(n2123) );
  NAND2X1 U1148 ( .A(\mem<20><1> ), .B(n104), .Y(n1443) );
  OAI21X1 U1149 ( .A(n103), .B(n1220), .C(n1443), .Y(n2122) );
  NAND2X1 U1150 ( .A(\mem<20><2> ), .B(n104), .Y(n1444) );
  OAI21X1 U1151 ( .A(n103), .B(n1222), .C(n1444), .Y(n2121) );
  NAND2X1 U1152 ( .A(\mem<20><3> ), .B(n104), .Y(n1445) );
  OAI21X1 U1153 ( .A(n103), .B(n1224), .C(n1445), .Y(n2120) );
  NAND2X1 U1154 ( .A(\mem<20><4> ), .B(n104), .Y(n1446) );
  OAI21X1 U1155 ( .A(n103), .B(n1226), .C(n1446), .Y(n2119) );
  NAND2X1 U1156 ( .A(\mem<20><5> ), .B(n104), .Y(n1447) );
  OAI21X1 U1157 ( .A(n103), .B(n1228), .C(n1447), .Y(n2118) );
  NAND2X1 U1158 ( .A(\mem<20><6> ), .B(n104), .Y(n1448) );
  OAI21X1 U1159 ( .A(n103), .B(n1230), .C(n1448), .Y(n2117) );
  NAND2X1 U1160 ( .A(\mem<20><7> ), .B(n104), .Y(n1449) );
  OAI21X1 U1161 ( .A(n103), .B(n1232), .C(n1449), .Y(n2116) );
  NAND2X1 U1162 ( .A(\mem<20><8> ), .B(n104), .Y(n1450) );
  OAI21X1 U1163 ( .A(n103), .B(n1234), .C(n1450), .Y(n2115) );
  NAND2X1 U1164 ( .A(\mem<20><9> ), .B(n104), .Y(n1451) );
  OAI21X1 U1165 ( .A(n103), .B(n1236), .C(n1451), .Y(n2114) );
  NAND2X1 U1166 ( .A(\mem<20><10> ), .B(n104), .Y(n1452) );
  OAI21X1 U1167 ( .A(n103), .B(n1238), .C(n1452), .Y(n2113) );
  NAND2X1 U1168 ( .A(\mem<20><11> ), .B(n104), .Y(n1453) );
  OAI21X1 U1169 ( .A(n103), .B(n1240), .C(n1453), .Y(n2112) );
  NAND2X1 U1170 ( .A(\mem<20><12> ), .B(n104), .Y(n1454) );
  OAI21X1 U1171 ( .A(n103), .B(n1242), .C(n1454), .Y(n2111) );
  NAND2X1 U1172 ( .A(\mem<20><13> ), .B(n104), .Y(n1455) );
  OAI21X1 U1173 ( .A(n103), .B(n1244), .C(n1455), .Y(n2110) );
  NAND2X1 U1174 ( .A(\mem<20><14> ), .B(n104), .Y(n1456) );
  OAI21X1 U1175 ( .A(n103), .B(n1246), .C(n1456), .Y(n2109) );
  NAND2X1 U1177 ( .A(\mem<20><15> ), .B(n104), .Y(n1457) );
  OAI21X1 U1178 ( .A(n103), .B(n1248), .C(n1457), .Y(n2108) );
  NAND2X1 U1179 ( .A(\mem<19><0> ), .B(n107), .Y(n1458) );
  OAI21X1 U1180 ( .A(n106), .B(n1218), .C(n1458), .Y(n2107) );
  NAND2X1 U1181 ( .A(\mem<19><1> ), .B(n107), .Y(n1459) );
  OAI21X1 U1182 ( .A(n106), .B(n1220), .C(n1459), .Y(n2106) );
  NAND2X1 U1183 ( .A(\mem<19><2> ), .B(n107), .Y(n1460) );
  OAI21X1 U1184 ( .A(n106), .B(n1222), .C(n1460), .Y(n2105) );
  NAND2X1 U1185 ( .A(\mem<19><3> ), .B(n107), .Y(n1461) );
  OAI21X1 U1186 ( .A(n106), .B(n1224), .C(n1461), .Y(n2104) );
  NAND2X1 U1187 ( .A(\mem<19><4> ), .B(n107), .Y(n1462) );
  OAI21X1 U1188 ( .A(n106), .B(n1226), .C(n1462), .Y(n2103) );
  NAND2X1 U1189 ( .A(\mem<19><5> ), .B(n107), .Y(n1463) );
  OAI21X1 U1190 ( .A(n106), .B(n1228), .C(n1463), .Y(n2102) );
  NAND2X1 U1191 ( .A(\mem<19><6> ), .B(n107), .Y(n1464) );
  OAI21X1 U1192 ( .A(n106), .B(n1230), .C(n1464), .Y(n2101) );
  NAND2X1 U1193 ( .A(\mem<19><7> ), .B(n107), .Y(n1465) );
  OAI21X1 U1194 ( .A(n106), .B(n1232), .C(n1465), .Y(n2100) );
  NAND2X1 U1195 ( .A(\mem<19><8> ), .B(n107), .Y(n1466) );
  OAI21X1 U1196 ( .A(n106), .B(n1234), .C(n1466), .Y(n2099) );
  NAND2X1 U1197 ( .A(\mem<19><9> ), .B(n107), .Y(n1467) );
  OAI21X1 U1198 ( .A(n106), .B(n1236), .C(n1467), .Y(n2098) );
  NAND2X1 U1199 ( .A(\mem<19><10> ), .B(n107), .Y(n1468) );
  OAI21X1 U1200 ( .A(n106), .B(n1238), .C(n1468), .Y(n2097) );
  NAND2X1 U1201 ( .A(\mem<19><11> ), .B(n107), .Y(n1469) );
  OAI21X1 U1202 ( .A(n106), .B(n1240), .C(n1469), .Y(n2096) );
  NAND2X1 U1203 ( .A(\mem<19><12> ), .B(n107), .Y(n1470) );
  OAI21X1 U1204 ( .A(n106), .B(n1242), .C(n1470), .Y(n2095) );
  NAND2X1 U1205 ( .A(\mem<19><13> ), .B(n107), .Y(n1471) );
  OAI21X1 U1206 ( .A(n106), .B(n1244), .C(n1471), .Y(n2094) );
  NAND2X1 U1207 ( .A(\mem<19><14> ), .B(n107), .Y(n1472) );
  OAI21X1 U1208 ( .A(n106), .B(n1246), .C(n1472), .Y(n2093) );
  NAND2X1 U1209 ( .A(\mem<19><15> ), .B(n107), .Y(n1473) );
  OAI21X1 U1210 ( .A(n106), .B(n1248), .C(n1473), .Y(n2092) );
  NAND2X1 U1211 ( .A(\mem<18><0> ), .B(n110), .Y(n1474) );
  OAI21X1 U1212 ( .A(n109), .B(n1218), .C(n1474), .Y(n2091) );
  NAND2X1 U1213 ( .A(\mem<18><1> ), .B(n110), .Y(n1475) );
  OAI21X1 U1214 ( .A(n109), .B(n1220), .C(n1475), .Y(n2090) );
  NAND2X1 U1215 ( .A(\mem<18><2> ), .B(n110), .Y(n1476) );
  OAI21X1 U1216 ( .A(n109), .B(n1222), .C(n1476), .Y(n2089) );
  NAND2X1 U1217 ( .A(\mem<18><3> ), .B(n110), .Y(n1477) );
  OAI21X1 U1218 ( .A(n109), .B(n1224), .C(n1477), .Y(n2088) );
  NAND2X1 U1219 ( .A(\mem<18><4> ), .B(n110), .Y(n1478) );
  OAI21X1 U1220 ( .A(n109), .B(n1226), .C(n1478), .Y(n2087) );
  NAND2X1 U1221 ( .A(\mem<18><5> ), .B(n110), .Y(n1479) );
  OAI21X1 U1222 ( .A(n109), .B(n1228), .C(n1479), .Y(n2086) );
  NAND2X1 U1223 ( .A(\mem<18><6> ), .B(n110), .Y(n1480) );
  OAI21X1 U1224 ( .A(n109), .B(n1230), .C(n1480), .Y(n2085) );
  NAND2X1 U1225 ( .A(\mem<18><7> ), .B(n110), .Y(n1481) );
  OAI21X1 U1226 ( .A(n109), .B(n1232), .C(n1481), .Y(n2084) );
  NAND2X1 U1227 ( .A(\mem<18><8> ), .B(n110), .Y(n1482) );
  OAI21X1 U1228 ( .A(n109), .B(n1234), .C(n1482), .Y(n2083) );
  NAND2X1 U1229 ( .A(\mem<18><9> ), .B(n110), .Y(n1483) );
  OAI21X1 U1230 ( .A(n109), .B(n1236), .C(n1483), .Y(n2082) );
  NAND2X1 U1231 ( .A(\mem<18><10> ), .B(n110), .Y(n1484) );
  OAI21X1 U1232 ( .A(n109), .B(n1238), .C(n1484), .Y(n2081) );
  NAND2X1 U1233 ( .A(\mem<18><11> ), .B(n110), .Y(n1485) );
  OAI21X1 U1234 ( .A(n109), .B(n1240), .C(n1485), .Y(n2080) );
  NAND2X1 U1235 ( .A(\mem<18><12> ), .B(n110), .Y(n1486) );
  OAI21X1 U1236 ( .A(n109), .B(n1242), .C(n1486), .Y(n2079) );
  NAND2X1 U1237 ( .A(\mem<18><13> ), .B(n110), .Y(n1487) );
  OAI21X1 U1238 ( .A(n109), .B(n1244), .C(n1487), .Y(n2078) );
  NAND2X1 U1239 ( .A(\mem<18><14> ), .B(n110), .Y(n1488) );
  OAI21X1 U1240 ( .A(n109), .B(n1246), .C(n1488), .Y(n2077) );
  NAND2X1 U1241 ( .A(\mem<18><15> ), .B(n110), .Y(n1489) );
  OAI21X1 U1242 ( .A(n109), .B(n1248), .C(n1489), .Y(n2076) );
  NAND2X1 U1243 ( .A(\mem<17><0> ), .B(n113), .Y(n1490) );
  OAI21X1 U1244 ( .A(n112), .B(n1218), .C(n1490), .Y(n2075) );
  NAND2X1 U1245 ( .A(\mem<17><1> ), .B(n113), .Y(n1491) );
  OAI21X1 U1246 ( .A(n112), .B(n1220), .C(n1491), .Y(n2074) );
  NAND2X1 U1247 ( .A(\mem<17><2> ), .B(n113), .Y(n1492) );
  OAI21X1 U1248 ( .A(n112), .B(n1222), .C(n1492), .Y(n2073) );
  NAND2X1 U1249 ( .A(\mem<17><3> ), .B(n113), .Y(n1493) );
  OAI21X1 U1250 ( .A(n112), .B(n1224), .C(n1493), .Y(n2072) );
  NAND2X1 U1251 ( .A(\mem<17><4> ), .B(n113), .Y(n1494) );
  OAI21X1 U1252 ( .A(n112), .B(n1226), .C(n1494), .Y(n2071) );
  NAND2X1 U1253 ( .A(\mem<17><5> ), .B(n113), .Y(n1495) );
  OAI21X1 U1254 ( .A(n112), .B(n1228), .C(n1495), .Y(n2070) );
  NAND2X1 U1255 ( .A(\mem<17><6> ), .B(n113), .Y(n1496) );
  OAI21X1 U1256 ( .A(n112), .B(n1230), .C(n1496), .Y(n2069) );
  NAND2X1 U1257 ( .A(\mem<17><7> ), .B(n113), .Y(n1497) );
  OAI21X1 U1258 ( .A(n112), .B(n1232), .C(n1497), .Y(n2068) );
  NAND2X1 U1259 ( .A(\mem<17><8> ), .B(n113), .Y(n1498) );
  OAI21X1 U1260 ( .A(n112), .B(n1234), .C(n1498), .Y(n2067) );
  NAND2X1 U1261 ( .A(\mem<17><9> ), .B(n113), .Y(n1499) );
  OAI21X1 U1262 ( .A(n112), .B(n1236), .C(n1499), .Y(n2066) );
  NAND2X1 U1263 ( .A(\mem<17><10> ), .B(n113), .Y(n1500) );
  OAI21X1 U1264 ( .A(n112), .B(n1238), .C(n1500), .Y(n2065) );
  NAND2X1 U1265 ( .A(\mem<17><11> ), .B(n113), .Y(n1501) );
  OAI21X1 U1266 ( .A(n112), .B(n1240), .C(n1501), .Y(n2064) );
  NAND2X1 U1267 ( .A(\mem<17><12> ), .B(n113), .Y(n1502) );
  OAI21X1 U1268 ( .A(n112), .B(n1242), .C(n1502), .Y(n2063) );
  NAND2X1 U1269 ( .A(\mem<17><13> ), .B(n113), .Y(n1503) );
  OAI21X1 U1270 ( .A(n112), .B(n1244), .C(n1503), .Y(n2062) );
  NAND2X1 U1271 ( .A(\mem<17><14> ), .B(n113), .Y(n1504) );
  OAI21X1 U1272 ( .A(n112), .B(n1246), .C(n1504), .Y(n2061) );
  NAND2X1 U1273 ( .A(\mem<17><15> ), .B(n113), .Y(n1505) );
  OAI21X1 U1274 ( .A(n112), .B(n1248), .C(n1505), .Y(n2060) );
  NAND2X1 U1275 ( .A(\mem<16><0> ), .B(n114), .Y(n1506) );
  OAI21X1 U1276 ( .A(n1209), .B(n1218), .C(n1506), .Y(n2059) );
  NAND2X1 U1277 ( .A(\mem<16><1> ), .B(n114), .Y(n1507) );
  OAI21X1 U1278 ( .A(n1209), .B(n1220), .C(n1507), .Y(n2058) );
  NAND2X1 U1279 ( .A(\mem<16><2> ), .B(n114), .Y(n1508) );
  OAI21X1 U1280 ( .A(n1209), .B(n1222), .C(n1508), .Y(n2057) );
  NAND2X1 U1281 ( .A(\mem<16><3> ), .B(n114), .Y(n1509) );
  OAI21X1 U1282 ( .A(n1209), .B(n1224), .C(n1509), .Y(n2056) );
  NAND2X1 U1283 ( .A(\mem<16><4> ), .B(n114), .Y(n1510) );
  OAI21X1 U1284 ( .A(n1209), .B(n1226), .C(n1510), .Y(n2055) );
  NAND2X1 U1285 ( .A(\mem<16><5> ), .B(n114), .Y(n1511) );
  OAI21X1 U1286 ( .A(n1209), .B(n1228), .C(n1511), .Y(n2054) );
  NAND2X1 U1287 ( .A(\mem<16><6> ), .B(n114), .Y(n1512) );
  OAI21X1 U1288 ( .A(n1209), .B(n1230), .C(n1512), .Y(n2053) );
  NAND2X1 U1289 ( .A(\mem<16><7> ), .B(n114), .Y(n1513) );
  OAI21X1 U1290 ( .A(n1209), .B(n1232), .C(n1513), .Y(n2052) );
  NAND2X1 U1291 ( .A(\mem<16><8> ), .B(n114), .Y(n1514) );
  OAI21X1 U1292 ( .A(n1209), .B(n1234), .C(n1514), .Y(n2051) );
  NAND2X1 U1293 ( .A(\mem<16><9> ), .B(n114), .Y(n1515) );
  OAI21X1 U1294 ( .A(n1209), .B(n1236), .C(n1515), .Y(n2050) );
  NAND2X1 U1295 ( .A(\mem<16><10> ), .B(n114), .Y(n1516) );
  OAI21X1 U1296 ( .A(n1209), .B(n1238), .C(n1516), .Y(n2049) );
  NAND2X1 U1297 ( .A(\mem<16><11> ), .B(n114), .Y(n1517) );
  OAI21X1 U1298 ( .A(n1209), .B(n1240), .C(n1517), .Y(n2048) );
  NAND2X1 U1299 ( .A(\mem<16><12> ), .B(n114), .Y(n1518) );
  OAI21X1 U1300 ( .A(n1209), .B(n1242), .C(n1518), .Y(n2047) );
  NAND2X1 U1301 ( .A(\mem<16><13> ), .B(n114), .Y(n1519) );
  OAI21X1 U1302 ( .A(n1209), .B(n1244), .C(n1519), .Y(n2046) );
  NAND2X1 U1303 ( .A(\mem<16><14> ), .B(n114), .Y(n1520) );
  OAI21X1 U1304 ( .A(n1209), .B(n1246), .C(n1520), .Y(n2045) );
  NAND2X1 U1305 ( .A(\mem<16><15> ), .B(n114), .Y(n1521) );
  OAI21X1 U1306 ( .A(n1209), .B(n1248), .C(n1521), .Y(n2044) );
  NAND3X1 U1307 ( .A(n1170), .B(n2300), .C(n1258), .Y(n1522) );
  NAND2X1 U1308 ( .A(\mem<15><0> ), .B(n117), .Y(n1523) );
  OAI21X1 U1309 ( .A(n116), .B(n1218), .C(n1523), .Y(n2043) );
  NAND2X1 U1310 ( .A(\mem<15><1> ), .B(n117), .Y(n1524) );
  OAI21X1 U1311 ( .A(n116), .B(n1220), .C(n1524), .Y(n2042) );
  NAND2X1 U1312 ( .A(\mem<15><2> ), .B(n117), .Y(n1525) );
  OAI21X1 U1313 ( .A(n116), .B(n1222), .C(n1525), .Y(n2041) );
  NAND2X1 U1314 ( .A(\mem<15><3> ), .B(n117), .Y(n1526) );
  OAI21X1 U1315 ( .A(n116), .B(n1224), .C(n1526), .Y(n2040) );
  NAND2X1 U1316 ( .A(\mem<15><4> ), .B(n117), .Y(n1527) );
  OAI21X1 U1317 ( .A(n116), .B(n1226), .C(n1527), .Y(n2039) );
  NAND2X1 U1318 ( .A(\mem<15><5> ), .B(n117), .Y(n1528) );
  OAI21X1 U1319 ( .A(n116), .B(n1228), .C(n1528), .Y(n2038) );
  NAND2X1 U1320 ( .A(\mem<15><6> ), .B(n117), .Y(n1529) );
  OAI21X1 U1321 ( .A(n116), .B(n1230), .C(n1529), .Y(n2037) );
  NAND2X1 U1322 ( .A(\mem<15><7> ), .B(n117), .Y(n1530) );
  OAI21X1 U1323 ( .A(n116), .B(n1232), .C(n1530), .Y(n2036) );
  NAND2X1 U1324 ( .A(\mem<15><8> ), .B(n117), .Y(n1531) );
  OAI21X1 U1325 ( .A(n116), .B(n1234), .C(n1531), .Y(n2035) );
  NAND2X1 U1326 ( .A(\mem<15><9> ), .B(n117), .Y(n1532) );
  OAI21X1 U1327 ( .A(n116), .B(n1236), .C(n1532), .Y(n2034) );
  NAND2X1 U1328 ( .A(\mem<15><10> ), .B(n117), .Y(n1533) );
  OAI21X1 U1329 ( .A(n116), .B(n1238), .C(n1533), .Y(n2033) );
  NAND2X1 U1330 ( .A(\mem<15><11> ), .B(n117), .Y(n1534) );
  OAI21X1 U1331 ( .A(n116), .B(n1240), .C(n1534), .Y(n2032) );
  NAND2X1 U1332 ( .A(\mem<15><12> ), .B(n117), .Y(n1535) );
  OAI21X1 U1333 ( .A(n116), .B(n1242), .C(n1535), .Y(n2031) );
  NAND2X1 U1334 ( .A(\mem<15><13> ), .B(n117), .Y(n1536) );
  OAI21X1 U1335 ( .A(n116), .B(n1244), .C(n1536), .Y(n2030) );
  NAND2X1 U1336 ( .A(\mem<15><14> ), .B(n117), .Y(n1537) );
  OAI21X1 U1337 ( .A(n116), .B(n1246), .C(n1537), .Y(n2029) );
  NAND2X1 U1338 ( .A(\mem<15><15> ), .B(n117), .Y(n1538) );
  OAI21X1 U1339 ( .A(n116), .B(n1248), .C(n1538), .Y(n2028) );
  NAND2X1 U1340 ( .A(\mem<14><0> ), .B(n120), .Y(n1539) );
  OAI21X1 U1341 ( .A(n119), .B(n1218), .C(n1539), .Y(n2027) );
  NAND2X1 U1342 ( .A(\mem<14><1> ), .B(n120), .Y(n1540) );
  OAI21X1 U1343 ( .A(n119), .B(n1220), .C(n1540), .Y(n2026) );
  NAND2X1 U1344 ( .A(\mem<14><2> ), .B(n120), .Y(n1541) );
  OAI21X1 U1345 ( .A(n119), .B(n1222), .C(n1541), .Y(n2025) );
  NAND2X1 U1346 ( .A(\mem<14><3> ), .B(n120), .Y(n1542) );
  OAI21X1 U1347 ( .A(n119), .B(n1224), .C(n1542), .Y(n2024) );
  NAND2X1 U1348 ( .A(\mem<14><4> ), .B(n120), .Y(n1543) );
  OAI21X1 U1349 ( .A(n119), .B(n1226), .C(n1543), .Y(n2023) );
  NAND2X1 U1350 ( .A(\mem<14><5> ), .B(n120), .Y(n1544) );
  OAI21X1 U1351 ( .A(n119), .B(n1228), .C(n1544), .Y(n2022) );
  NAND2X1 U1352 ( .A(\mem<14><6> ), .B(n120), .Y(n1545) );
  OAI21X1 U1353 ( .A(n119), .B(n1230), .C(n1545), .Y(n2021) );
  NAND2X1 U1354 ( .A(\mem<14><7> ), .B(n120), .Y(n1546) );
  OAI21X1 U1355 ( .A(n119), .B(n1232), .C(n1546), .Y(n2020) );
  NAND2X1 U1356 ( .A(\mem<14><8> ), .B(n120), .Y(n1547) );
  OAI21X1 U1357 ( .A(n119), .B(n1234), .C(n1547), .Y(n2019) );
  NAND2X1 U1358 ( .A(\mem<14><9> ), .B(n120), .Y(n1548) );
  OAI21X1 U1359 ( .A(n119), .B(n1236), .C(n1548), .Y(n2018) );
  NAND2X1 U1360 ( .A(\mem<14><10> ), .B(n120), .Y(n1549) );
  OAI21X1 U1361 ( .A(n119), .B(n1238), .C(n1549), .Y(n2017) );
  NAND2X1 U1362 ( .A(\mem<14><11> ), .B(n120), .Y(n1550) );
  OAI21X1 U1363 ( .A(n119), .B(n1240), .C(n1550), .Y(n2016) );
  NAND2X1 U1364 ( .A(\mem<14><12> ), .B(n120), .Y(n1551) );
  OAI21X1 U1365 ( .A(n119), .B(n1242), .C(n1551), .Y(n2015) );
  NAND2X1 U1366 ( .A(\mem<14><13> ), .B(n120), .Y(n1552) );
  OAI21X1 U1367 ( .A(n119), .B(n1244), .C(n1552), .Y(n2014) );
  NAND2X1 U1368 ( .A(\mem<14><14> ), .B(n120), .Y(n1553) );
  OAI21X1 U1369 ( .A(n119), .B(n1246), .C(n1553), .Y(n2013) );
  NAND2X1 U1370 ( .A(\mem<14><15> ), .B(n120), .Y(n1554) );
  OAI21X1 U1371 ( .A(n119), .B(n1248), .C(n1554), .Y(n2012) );
  NAND2X1 U1372 ( .A(\mem<13><0> ), .B(n123), .Y(n1555) );
  OAI21X1 U1373 ( .A(n122), .B(n1218), .C(n1555), .Y(n2011) );
  NAND2X1 U1374 ( .A(\mem<13><1> ), .B(n123), .Y(n1556) );
  OAI21X1 U1375 ( .A(n122), .B(n1220), .C(n1556), .Y(n2010) );
  NAND2X1 U1376 ( .A(\mem<13><2> ), .B(n123), .Y(n1557) );
  OAI21X1 U1377 ( .A(n122), .B(n1222), .C(n1557), .Y(n2009) );
  NAND2X1 U1378 ( .A(\mem<13><3> ), .B(n123), .Y(n1558) );
  OAI21X1 U1379 ( .A(n122), .B(n1224), .C(n1558), .Y(n2008) );
  NAND2X1 U1380 ( .A(\mem<13><4> ), .B(n123), .Y(n1559) );
  OAI21X1 U1381 ( .A(n122), .B(n1226), .C(n1559), .Y(n2007) );
  NAND2X1 U1382 ( .A(\mem<13><5> ), .B(n123), .Y(n1560) );
  OAI21X1 U1383 ( .A(n122), .B(n1228), .C(n1560), .Y(n2006) );
  NAND2X1 U1384 ( .A(\mem<13><6> ), .B(n123), .Y(n1561) );
  OAI21X1 U1385 ( .A(n122), .B(n1230), .C(n1561), .Y(n2005) );
  NAND2X1 U1386 ( .A(\mem<13><7> ), .B(n123), .Y(n1562) );
  OAI21X1 U1387 ( .A(n122), .B(n1232), .C(n1562), .Y(n2004) );
  NAND2X1 U1388 ( .A(\mem<13><8> ), .B(n123), .Y(n1563) );
  OAI21X1 U1389 ( .A(n122), .B(n1234), .C(n1563), .Y(n2003) );
  NAND2X1 U1390 ( .A(\mem<13><9> ), .B(n123), .Y(n1564) );
  OAI21X1 U1391 ( .A(n122), .B(n1236), .C(n1564), .Y(n2002) );
  NAND2X1 U1392 ( .A(\mem<13><10> ), .B(n123), .Y(n1565) );
  OAI21X1 U1393 ( .A(n122), .B(n1238), .C(n1565), .Y(n2001) );
  NAND2X1 U1394 ( .A(\mem<13><11> ), .B(n123), .Y(n1566) );
  OAI21X1 U1395 ( .A(n122), .B(n1240), .C(n1566), .Y(n2000) );
  NAND2X1 U1396 ( .A(\mem<13><12> ), .B(n123), .Y(n1567) );
  OAI21X1 U1397 ( .A(n122), .B(n1242), .C(n1567), .Y(n1999) );
  NAND2X1 U1398 ( .A(\mem<13><13> ), .B(n123), .Y(n1568) );
  OAI21X1 U1399 ( .A(n122), .B(n1244), .C(n1568), .Y(n1998) );
  NAND2X1 U1400 ( .A(\mem<13><14> ), .B(n123), .Y(n1569) );
  OAI21X1 U1401 ( .A(n122), .B(n1246), .C(n1569), .Y(n1997) );
  NAND2X1 U1402 ( .A(\mem<13><15> ), .B(n123), .Y(n1570) );
  OAI21X1 U1403 ( .A(n122), .B(n1248), .C(n1570), .Y(n1996) );
  NAND2X1 U1404 ( .A(\mem<12><0> ), .B(n126), .Y(n1571) );
  OAI21X1 U1405 ( .A(n125), .B(n1218), .C(n1571), .Y(n1995) );
  NAND2X1 U1406 ( .A(\mem<12><1> ), .B(n126), .Y(n1572) );
  OAI21X1 U1407 ( .A(n125), .B(n1220), .C(n1572), .Y(n1994) );
  NAND2X1 U1408 ( .A(\mem<12><2> ), .B(n126), .Y(n1573) );
  OAI21X1 U1409 ( .A(n125), .B(n1222), .C(n1573), .Y(n1993) );
  NAND2X1 U1410 ( .A(\mem<12><3> ), .B(n126), .Y(n1574) );
  OAI21X1 U1411 ( .A(n125), .B(n1224), .C(n1574), .Y(n1992) );
  NAND2X1 U1412 ( .A(\mem<12><4> ), .B(n126), .Y(n1575) );
  OAI21X1 U1413 ( .A(n125), .B(n1226), .C(n1575), .Y(n1991) );
  NAND2X1 U1414 ( .A(\mem<12><5> ), .B(n126), .Y(n1576) );
  OAI21X1 U1415 ( .A(n125), .B(n1228), .C(n1576), .Y(n1990) );
  NAND2X1 U1416 ( .A(\mem<12><6> ), .B(n126), .Y(n1577) );
  OAI21X1 U1417 ( .A(n125), .B(n1230), .C(n1577), .Y(n1989) );
  NAND2X1 U1418 ( .A(\mem<12><7> ), .B(n126), .Y(n1578) );
  OAI21X1 U1419 ( .A(n125), .B(n1232), .C(n1578), .Y(n1988) );
  NAND2X1 U1420 ( .A(\mem<12><8> ), .B(n126), .Y(n1579) );
  OAI21X1 U1421 ( .A(n125), .B(n1234), .C(n1579), .Y(n1987) );
  NAND2X1 U1422 ( .A(\mem<12><9> ), .B(n126), .Y(n1580) );
  OAI21X1 U1423 ( .A(n125), .B(n1236), .C(n1580), .Y(n1986) );
  NAND2X1 U1424 ( .A(\mem<12><10> ), .B(n126), .Y(n1581) );
  OAI21X1 U1425 ( .A(n125), .B(n1238), .C(n1581), .Y(n1985) );
  NAND2X1 U1426 ( .A(\mem<12><11> ), .B(n126), .Y(n1582) );
  OAI21X1 U1427 ( .A(n125), .B(n1240), .C(n1582), .Y(n1984) );
  NAND2X1 U1428 ( .A(\mem<12><12> ), .B(n126), .Y(n1583) );
  OAI21X1 U1429 ( .A(n125), .B(n1242), .C(n1583), .Y(n1983) );
  NAND2X1 U1430 ( .A(\mem<12><13> ), .B(n126), .Y(n1584) );
  OAI21X1 U1431 ( .A(n125), .B(n1244), .C(n1584), .Y(n1982) );
  NAND2X1 U1432 ( .A(\mem<12><14> ), .B(n126), .Y(n1585) );
  OAI21X1 U1433 ( .A(n125), .B(n1246), .C(n1585), .Y(n1981) );
  NAND2X1 U1434 ( .A(\mem<12><15> ), .B(n126), .Y(n1586) );
  OAI21X1 U1435 ( .A(n125), .B(n1248), .C(n1586), .Y(n1980) );
  NAND2X1 U1436 ( .A(\mem<11><0> ), .B(n129), .Y(n1587) );
  OAI21X1 U1437 ( .A(n128), .B(n1218), .C(n1587), .Y(n1979) );
  NAND2X1 U1438 ( .A(\mem<11><1> ), .B(n129), .Y(n1588) );
  OAI21X1 U1439 ( .A(n128), .B(n1219), .C(n1588), .Y(n1978) );
  NAND2X1 U1440 ( .A(\mem<11><2> ), .B(n129), .Y(n1589) );
  OAI21X1 U1441 ( .A(n128), .B(n1221), .C(n1589), .Y(n1977) );
  NAND2X1 U1442 ( .A(\mem<11><3> ), .B(n129), .Y(n1590) );
  OAI21X1 U1443 ( .A(n128), .B(n1223), .C(n1590), .Y(n1976) );
  NAND2X1 U1444 ( .A(\mem<11><4> ), .B(n129), .Y(n1591) );
  OAI21X1 U1445 ( .A(n128), .B(n1225), .C(n1591), .Y(n1975) );
  NAND2X1 U1446 ( .A(\mem<11><5> ), .B(n129), .Y(n1592) );
  OAI21X1 U1447 ( .A(n128), .B(n1227), .C(n1592), .Y(n1974) );
  NAND2X1 U1448 ( .A(\mem<11><6> ), .B(n129), .Y(n1593) );
  OAI21X1 U1449 ( .A(n128), .B(n1229), .C(n1593), .Y(n1973) );
  NAND2X1 U1450 ( .A(\mem<11><7> ), .B(n129), .Y(n1594) );
  OAI21X1 U1451 ( .A(n128), .B(n1231), .C(n1594), .Y(n1972) );
  NAND2X1 U1452 ( .A(\mem<11><8> ), .B(n129), .Y(n1595) );
  OAI21X1 U1453 ( .A(n128), .B(n1233), .C(n1595), .Y(n1971) );
  NAND2X1 U1454 ( .A(\mem<11><9> ), .B(n129), .Y(n1596) );
  OAI21X1 U1455 ( .A(n128), .B(n1235), .C(n1596), .Y(n1970) );
  NAND2X1 U1456 ( .A(\mem<11><10> ), .B(n129), .Y(n1597) );
  OAI21X1 U1457 ( .A(n128), .B(n1237), .C(n1597), .Y(n1969) );
  NAND2X1 U1458 ( .A(\mem<11><11> ), .B(n129), .Y(n1598) );
  OAI21X1 U1459 ( .A(n128), .B(n1239), .C(n1598), .Y(n1968) );
  NAND2X1 U1460 ( .A(\mem<11><12> ), .B(n129), .Y(n1599) );
  OAI21X1 U1461 ( .A(n128), .B(n1241), .C(n1599), .Y(n1967) );
  NAND2X1 U1462 ( .A(\mem<11><13> ), .B(n129), .Y(n1600) );
  OAI21X1 U1463 ( .A(n128), .B(n1243), .C(n1600), .Y(n1966) );
  NAND2X1 U1464 ( .A(\mem<11><14> ), .B(n129), .Y(n1601) );
  OAI21X1 U1465 ( .A(n128), .B(n1245), .C(n1601), .Y(n1965) );
  NAND2X1 U1466 ( .A(\mem<11><15> ), .B(n129), .Y(n1602) );
  OAI21X1 U1467 ( .A(n128), .B(n1247), .C(n1602), .Y(n1964) );
  NAND2X1 U1468 ( .A(\mem<10><0> ), .B(n132), .Y(n1603) );
  OAI21X1 U1469 ( .A(n131), .B(n1218), .C(n1603), .Y(n1963) );
  NAND2X1 U1470 ( .A(\mem<10><1> ), .B(n132), .Y(n1604) );
  OAI21X1 U1471 ( .A(n131), .B(n1219), .C(n1604), .Y(n1962) );
  NAND2X1 U1472 ( .A(\mem<10><2> ), .B(n132), .Y(n1605) );
  OAI21X1 U1473 ( .A(n131), .B(n1221), .C(n1605), .Y(n1961) );
  NAND2X1 U1474 ( .A(\mem<10><3> ), .B(n132), .Y(n1606) );
  OAI21X1 U1475 ( .A(n131), .B(n1223), .C(n1606), .Y(n1960) );
  NAND2X1 U1476 ( .A(\mem<10><4> ), .B(n132), .Y(n1607) );
  OAI21X1 U1477 ( .A(n131), .B(n1225), .C(n1607), .Y(n1959) );
  NAND2X1 U1478 ( .A(\mem<10><5> ), .B(n132), .Y(n1608) );
  OAI21X1 U1479 ( .A(n131), .B(n1227), .C(n1608), .Y(n1958) );
  NAND2X1 U1480 ( .A(\mem<10><6> ), .B(n132), .Y(n1609) );
  OAI21X1 U1481 ( .A(n131), .B(n1229), .C(n1609), .Y(n1957) );
  NAND2X1 U1482 ( .A(\mem<10><7> ), .B(n132), .Y(n1610) );
  OAI21X1 U1483 ( .A(n131), .B(n1231), .C(n1610), .Y(n1956) );
  NAND2X1 U1484 ( .A(\mem<10><8> ), .B(n132), .Y(n1611) );
  OAI21X1 U1485 ( .A(n131), .B(n1233), .C(n1611), .Y(n1955) );
  NAND2X1 U1486 ( .A(\mem<10><9> ), .B(n132), .Y(n1612) );
  OAI21X1 U1487 ( .A(n131), .B(n1235), .C(n1612), .Y(n1954) );
  NAND2X1 U1488 ( .A(\mem<10><10> ), .B(n132), .Y(n1613) );
  OAI21X1 U1489 ( .A(n131), .B(n1237), .C(n1613), .Y(n1953) );
  NAND2X1 U1490 ( .A(\mem<10><11> ), .B(n132), .Y(n1614) );
  OAI21X1 U1491 ( .A(n131), .B(n1239), .C(n1614), .Y(n1952) );
  NAND2X1 U1492 ( .A(\mem<10><12> ), .B(n132), .Y(n1615) );
  OAI21X1 U1493 ( .A(n131), .B(n1241), .C(n1615), .Y(n1951) );
  NAND2X1 U1494 ( .A(\mem<10><13> ), .B(n132), .Y(n1616) );
  OAI21X1 U1495 ( .A(n131), .B(n1243), .C(n1616), .Y(n1950) );
  NAND2X1 U1496 ( .A(\mem<10><14> ), .B(n132), .Y(n1617) );
  OAI21X1 U1497 ( .A(n131), .B(n1245), .C(n1617), .Y(n1949) );
  NAND2X1 U1498 ( .A(\mem<10><15> ), .B(n132), .Y(n1618) );
  OAI21X1 U1499 ( .A(n131), .B(n1247), .C(n1618), .Y(n1948) );
  NAND2X1 U1500 ( .A(\mem<9><0> ), .B(n135), .Y(n1619) );
  OAI21X1 U1501 ( .A(n134), .B(n1218), .C(n1619), .Y(n1947) );
  NAND2X1 U1502 ( .A(\mem<9><1> ), .B(n135), .Y(n1620) );
  OAI21X1 U1503 ( .A(n134), .B(n1219), .C(n1620), .Y(n1946) );
  NAND2X1 U1504 ( .A(\mem<9><2> ), .B(n135), .Y(n1621) );
  OAI21X1 U1505 ( .A(n134), .B(n1221), .C(n1621), .Y(n1945) );
  NAND2X1 U1506 ( .A(\mem<9><3> ), .B(n135), .Y(n1622) );
  OAI21X1 U1507 ( .A(n134), .B(n1223), .C(n1622), .Y(n1944) );
  NAND2X1 U1508 ( .A(\mem<9><4> ), .B(n135), .Y(n1623) );
  OAI21X1 U1509 ( .A(n134), .B(n1225), .C(n1623), .Y(n1943) );
  NAND2X1 U1510 ( .A(\mem<9><5> ), .B(n135), .Y(n1624) );
  OAI21X1 U1511 ( .A(n134), .B(n1227), .C(n1624), .Y(n1942) );
  NAND2X1 U1512 ( .A(\mem<9><6> ), .B(n135), .Y(n1625) );
  OAI21X1 U1513 ( .A(n134), .B(n1229), .C(n1625), .Y(n1941) );
  NAND2X1 U1514 ( .A(\mem<9><7> ), .B(n135), .Y(n1626) );
  OAI21X1 U1515 ( .A(n134), .B(n1231), .C(n1626), .Y(n1940) );
  NAND2X1 U1516 ( .A(\mem<9><8> ), .B(n135), .Y(n1627) );
  OAI21X1 U1517 ( .A(n134), .B(n1233), .C(n1627), .Y(n1939) );
  NAND2X1 U1518 ( .A(\mem<9><9> ), .B(n135), .Y(n1628) );
  OAI21X1 U1519 ( .A(n134), .B(n1235), .C(n1628), .Y(n1938) );
  NAND2X1 U1520 ( .A(\mem<9><10> ), .B(n135), .Y(n1629) );
  OAI21X1 U1521 ( .A(n134), .B(n1237), .C(n1629), .Y(n1937) );
  NAND2X1 U1522 ( .A(\mem<9><11> ), .B(n135), .Y(n1630) );
  OAI21X1 U1523 ( .A(n134), .B(n1239), .C(n1630), .Y(n1936) );
  NAND2X1 U1524 ( .A(\mem<9><12> ), .B(n135), .Y(n1631) );
  OAI21X1 U1525 ( .A(n134), .B(n1241), .C(n1631), .Y(n1935) );
  NAND2X1 U1526 ( .A(\mem<9><13> ), .B(n135), .Y(n1632) );
  OAI21X1 U1527 ( .A(n134), .B(n1243), .C(n1632), .Y(n1934) );
  NAND2X1 U1528 ( .A(\mem<9><14> ), .B(n135), .Y(n1633) );
  OAI21X1 U1529 ( .A(n134), .B(n1245), .C(n1633), .Y(n1933) );
  NAND2X1 U1530 ( .A(\mem<9><15> ), .B(n135), .Y(n1634) );
  OAI21X1 U1531 ( .A(n134), .B(n1247), .C(n1634), .Y(n1932) );
  NAND2X1 U1532 ( .A(\mem<8><0> ), .B(n136), .Y(n1636) );
  OAI21X1 U1533 ( .A(n1210), .B(n1218), .C(n1636), .Y(n1931) );
  NAND2X1 U1534 ( .A(\mem<8><1> ), .B(n136), .Y(n1637) );
  OAI21X1 U1535 ( .A(n1210), .B(n1219), .C(n1637), .Y(n1930) );
  NAND2X1 U1536 ( .A(\mem<8><2> ), .B(n136), .Y(n1638) );
  OAI21X1 U1537 ( .A(n1210), .B(n1221), .C(n1638), .Y(n1929) );
  NAND2X1 U1538 ( .A(\mem<8><3> ), .B(n136), .Y(n1639) );
  OAI21X1 U1539 ( .A(n1210), .B(n1223), .C(n1639), .Y(n1928) );
  NAND2X1 U1540 ( .A(\mem<8><4> ), .B(n136), .Y(n1640) );
  OAI21X1 U1541 ( .A(n1210), .B(n1225), .C(n1640), .Y(n1927) );
  NAND2X1 U1542 ( .A(\mem<8><5> ), .B(n136), .Y(n1641) );
  OAI21X1 U1543 ( .A(n1210), .B(n1227), .C(n1641), .Y(n1926) );
  NAND2X1 U1544 ( .A(\mem<8><6> ), .B(n136), .Y(n1642) );
  OAI21X1 U1545 ( .A(n1210), .B(n1229), .C(n1642), .Y(n1925) );
  NAND2X1 U1546 ( .A(\mem<8><7> ), .B(n136), .Y(n1643) );
  OAI21X1 U1547 ( .A(n1210), .B(n1231), .C(n1643), .Y(n1924) );
  NAND2X1 U1548 ( .A(\mem<8><8> ), .B(n136), .Y(n1644) );
  OAI21X1 U1549 ( .A(n1210), .B(n1233), .C(n1644), .Y(n1923) );
  NAND2X1 U1550 ( .A(\mem<8><9> ), .B(n136), .Y(n1645) );
  OAI21X1 U1551 ( .A(n1210), .B(n1235), .C(n1645), .Y(n1922) );
  NAND2X1 U1552 ( .A(\mem<8><10> ), .B(n136), .Y(n1646) );
  OAI21X1 U1553 ( .A(n1210), .B(n1237), .C(n1646), .Y(n1921) );
  NAND2X1 U1554 ( .A(\mem<8><11> ), .B(n136), .Y(n1647) );
  OAI21X1 U1555 ( .A(n1210), .B(n1239), .C(n1647), .Y(n1920) );
  NAND2X1 U1556 ( .A(\mem<8><12> ), .B(n136), .Y(n1648) );
  OAI21X1 U1557 ( .A(n1210), .B(n1241), .C(n1648), .Y(n1919) );
  NAND2X1 U1558 ( .A(\mem<8><13> ), .B(n136), .Y(n1649) );
  OAI21X1 U1559 ( .A(n1210), .B(n1243), .C(n1649), .Y(n1918) );
  NAND2X1 U1560 ( .A(\mem<8><14> ), .B(n136), .Y(n1650) );
  OAI21X1 U1561 ( .A(n1210), .B(n1245), .C(n1650), .Y(n1917) );
  NAND2X1 U1562 ( .A(\mem<8><15> ), .B(n136), .Y(n1651) );
  OAI21X1 U1563 ( .A(n1210), .B(n1247), .C(n1651), .Y(n1916) );
  NAND3X1 U1564 ( .A(n1256), .B(n2300), .C(n1258), .Y(n1652) );
  NAND2X1 U1565 ( .A(\mem<7><0> ), .B(n139), .Y(n1653) );
  OAI21X1 U1566 ( .A(n138), .B(n1217), .C(n1653), .Y(n1915) );
  NAND2X1 U1567 ( .A(\mem<7><1> ), .B(n139), .Y(n1654) );
  OAI21X1 U1568 ( .A(n138), .B(n1219), .C(n1654), .Y(n1914) );
  NAND2X1 U1569 ( .A(\mem<7><2> ), .B(n139), .Y(n1655) );
  OAI21X1 U1570 ( .A(n138), .B(n1221), .C(n1655), .Y(n1913) );
  NAND2X1 U1571 ( .A(\mem<7><3> ), .B(n139), .Y(n1656) );
  OAI21X1 U1572 ( .A(n138), .B(n1223), .C(n1656), .Y(n1912) );
  NAND2X1 U1573 ( .A(\mem<7><4> ), .B(n139), .Y(n1657) );
  OAI21X1 U1574 ( .A(n138), .B(n1225), .C(n1657), .Y(n1911) );
  NAND2X1 U1575 ( .A(\mem<7><5> ), .B(n139), .Y(n1658) );
  OAI21X1 U1576 ( .A(n138), .B(n1227), .C(n1658), .Y(n1910) );
  NAND2X1 U1577 ( .A(\mem<7><6> ), .B(n139), .Y(n1659) );
  OAI21X1 U1578 ( .A(n138), .B(n1229), .C(n1659), .Y(n1909) );
  NAND2X1 U1579 ( .A(\mem<7><7> ), .B(n139), .Y(n1660) );
  OAI21X1 U1580 ( .A(n138), .B(n1231), .C(n1660), .Y(n1908) );
  NAND2X1 U1581 ( .A(\mem<7><8> ), .B(n139), .Y(n1661) );
  OAI21X1 U1582 ( .A(n138), .B(n1233), .C(n1661), .Y(n1907) );
  NAND2X1 U1583 ( .A(\mem<7><9> ), .B(n139), .Y(n1662) );
  OAI21X1 U1584 ( .A(n138), .B(n1235), .C(n1662), .Y(n1906) );
  NAND2X1 U1585 ( .A(\mem<7><10> ), .B(n139), .Y(n1663) );
  OAI21X1 U1586 ( .A(n138), .B(n1237), .C(n1663), .Y(n1905) );
  NAND2X1 U1587 ( .A(\mem<7><11> ), .B(n139), .Y(n1664) );
  OAI21X1 U1588 ( .A(n138), .B(n1239), .C(n1664), .Y(n1904) );
  NAND2X1 U1589 ( .A(\mem<7><12> ), .B(n139), .Y(n1665) );
  OAI21X1 U1590 ( .A(n138), .B(n1241), .C(n1665), .Y(n1903) );
  NAND2X1 U1591 ( .A(\mem<7><13> ), .B(n139), .Y(n1666) );
  OAI21X1 U1592 ( .A(n138), .B(n1243), .C(n1666), .Y(n1902) );
  NAND2X1 U1593 ( .A(\mem<7><14> ), .B(n139), .Y(n1667) );
  OAI21X1 U1594 ( .A(n138), .B(n1245), .C(n1667), .Y(n1901) );
  NAND2X1 U1595 ( .A(\mem<7><15> ), .B(n139), .Y(n1668) );
  OAI21X1 U1596 ( .A(n138), .B(n1247), .C(n1668), .Y(n1900) );
  NAND2X1 U1597 ( .A(\mem<6><0> ), .B(n142), .Y(n1669) );
  OAI21X1 U1598 ( .A(n141), .B(n1218), .C(n1669), .Y(n1899) );
  NAND2X1 U1599 ( .A(\mem<6><1> ), .B(n142), .Y(n1670) );
  OAI21X1 U1600 ( .A(n141), .B(n1219), .C(n1670), .Y(n1898) );
  NAND2X1 U1601 ( .A(\mem<6><2> ), .B(n142), .Y(n1671) );
  OAI21X1 U1602 ( .A(n141), .B(n1221), .C(n1671), .Y(n1897) );
  NAND2X1 U1603 ( .A(\mem<6><3> ), .B(n142), .Y(n1672) );
  OAI21X1 U1604 ( .A(n141), .B(n1223), .C(n1672), .Y(n1896) );
  NAND2X1 U1605 ( .A(\mem<6><4> ), .B(n142), .Y(n1673) );
  OAI21X1 U1606 ( .A(n141), .B(n1225), .C(n1673), .Y(n1895) );
  NAND2X1 U1607 ( .A(\mem<6><5> ), .B(n142), .Y(n1674) );
  OAI21X1 U1608 ( .A(n141), .B(n1227), .C(n1674), .Y(n1894) );
  NAND2X1 U1609 ( .A(\mem<6><6> ), .B(n142), .Y(n1675) );
  OAI21X1 U1610 ( .A(n141), .B(n1229), .C(n1675), .Y(n1893) );
  NAND2X1 U1611 ( .A(\mem<6><7> ), .B(n142), .Y(n1676) );
  OAI21X1 U1612 ( .A(n141), .B(n1231), .C(n1676), .Y(n1892) );
  NAND2X1 U1613 ( .A(\mem<6><8> ), .B(n142), .Y(n1677) );
  OAI21X1 U1614 ( .A(n141), .B(n1233), .C(n1677), .Y(n1891) );
  NAND2X1 U1615 ( .A(\mem<6><9> ), .B(n142), .Y(n1678) );
  OAI21X1 U1616 ( .A(n141), .B(n1235), .C(n1678), .Y(n1890) );
  NAND2X1 U1617 ( .A(\mem<6><10> ), .B(n142), .Y(n1679) );
  OAI21X1 U1618 ( .A(n141), .B(n1237), .C(n1679), .Y(n1889) );
  NAND2X1 U1619 ( .A(\mem<6><11> ), .B(n142), .Y(n1680) );
  OAI21X1 U1620 ( .A(n141), .B(n1239), .C(n1680), .Y(n1888) );
  NAND2X1 U1621 ( .A(\mem<6><12> ), .B(n142), .Y(n1681) );
  OAI21X1 U1622 ( .A(n141), .B(n1241), .C(n1681), .Y(n1887) );
  NAND2X1 U1623 ( .A(\mem<6><13> ), .B(n142), .Y(n1682) );
  OAI21X1 U1624 ( .A(n141), .B(n1243), .C(n1682), .Y(n1886) );
  NAND2X1 U1625 ( .A(\mem<6><14> ), .B(n142), .Y(n1683) );
  OAI21X1 U1626 ( .A(n141), .B(n1245), .C(n1683), .Y(n1885) );
  NAND2X1 U1627 ( .A(\mem<6><15> ), .B(n142), .Y(n1684) );
  OAI21X1 U1628 ( .A(n141), .B(n1247), .C(n1684), .Y(n1884) );
  NAND2X1 U1629 ( .A(\mem<5><0> ), .B(n145), .Y(n1686) );
  OAI21X1 U1630 ( .A(n144), .B(n1217), .C(n1686), .Y(n1883) );
  NAND2X1 U1631 ( .A(\mem<5><1> ), .B(n145), .Y(n1687) );
  OAI21X1 U1632 ( .A(n144), .B(n1219), .C(n1687), .Y(n1882) );
  NAND2X1 U1633 ( .A(\mem<5><2> ), .B(n145), .Y(n1688) );
  OAI21X1 U1634 ( .A(n144), .B(n1221), .C(n1688), .Y(n1881) );
  NAND2X1 U1635 ( .A(\mem<5><3> ), .B(n145), .Y(n1689) );
  OAI21X1 U1636 ( .A(n144), .B(n1223), .C(n1689), .Y(n1880) );
  NAND2X1 U1637 ( .A(\mem<5><4> ), .B(n145), .Y(n1690) );
  OAI21X1 U1638 ( .A(n144), .B(n1225), .C(n1690), .Y(n1879) );
  NAND2X1 U1639 ( .A(\mem<5><5> ), .B(n145), .Y(n1691) );
  OAI21X1 U1640 ( .A(n144), .B(n1227), .C(n1691), .Y(n1878) );
  NAND2X1 U1641 ( .A(\mem<5><6> ), .B(n145), .Y(n1692) );
  OAI21X1 U1642 ( .A(n144), .B(n1229), .C(n1692), .Y(n1877) );
  NAND2X1 U1643 ( .A(\mem<5><7> ), .B(n145), .Y(n1693) );
  OAI21X1 U1644 ( .A(n144), .B(n1231), .C(n1693), .Y(n1876) );
  NAND2X1 U1645 ( .A(\mem<5><8> ), .B(n145), .Y(n1694) );
  OAI21X1 U1646 ( .A(n144), .B(n1233), .C(n1694), .Y(n1875) );
  NAND2X1 U1647 ( .A(\mem<5><9> ), .B(n145), .Y(n1695) );
  OAI21X1 U1648 ( .A(n144), .B(n1235), .C(n1695), .Y(n1874) );
  NAND2X1 U1649 ( .A(\mem<5><10> ), .B(n145), .Y(n1696) );
  OAI21X1 U1650 ( .A(n144), .B(n1237), .C(n1696), .Y(n1873) );
  NAND2X1 U1651 ( .A(\mem<5><11> ), .B(n145), .Y(n1697) );
  OAI21X1 U1652 ( .A(n144), .B(n1239), .C(n1697), .Y(n1872) );
  NAND2X1 U1653 ( .A(\mem<5><12> ), .B(n145), .Y(n1698) );
  OAI21X1 U1654 ( .A(n144), .B(n1241), .C(n1698), .Y(n1871) );
  NAND2X1 U1655 ( .A(\mem<5><13> ), .B(n145), .Y(n1699) );
  OAI21X1 U1656 ( .A(n144), .B(n1243), .C(n1699), .Y(n1870) );
  NAND2X1 U1657 ( .A(\mem<5><14> ), .B(n145), .Y(n1700) );
  OAI21X1 U1658 ( .A(n144), .B(n1245), .C(n1700), .Y(n1869) );
  NAND2X1 U1659 ( .A(\mem<5><15> ), .B(n145), .Y(n1701) );
  OAI21X1 U1660 ( .A(n144), .B(n1247), .C(n1701), .Y(n1868) );
  NAND2X1 U1661 ( .A(\mem<4><0> ), .B(n148), .Y(n1703) );
  OAI21X1 U1662 ( .A(n147), .B(n1218), .C(n1703), .Y(n1867) );
  NAND2X1 U1663 ( .A(\mem<4><1> ), .B(n148), .Y(n1704) );
  OAI21X1 U1664 ( .A(n147), .B(n1219), .C(n1704), .Y(n1866) );
  NAND2X1 U1665 ( .A(\mem<4><2> ), .B(n148), .Y(n1705) );
  OAI21X1 U1666 ( .A(n147), .B(n1221), .C(n1705), .Y(n1865) );
  NAND2X1 U1667 ( .A(\mem<4><3> ), .B(n148), .Y(n1706) );
  OAI21X1 U1668 ( .A(n147), .B(n1223), .C(n1706), .Y(n1864) );
  NAND2X1 U1669 ( .A(\mem<4><4> ), .B(n148), .Y(n1707) );
  OAI21X1 U1670 ( .A(n147), .B(n1225), .C(n1707), .Y(n1863) );
  NAND2X1 U1671 ( .A(\mem<4><5> ), .B(n148), .Y(n1708) );
  OAI21X1 U1672 ( .A(n147), .B(n1227), .C(n1708), .Y(n1862) );
  NAND2X1 U1673 ( .A(\mem<4><6> ), .B(n148), .Y(n1709) );
  OAI21X1 U1674 ( .A(n147), .B(n1229), .C(n1709), .Y(n1861) );
  NAND2X1 U1675 ( .A(\mem<4><7> ), .B(n148), .Y(n1710) );
  OAI21X1 U1676 ( .A(n147), .B(n1231), .C(n1710), .Y(n1860) );
  NAND2X1 U1677 ( .A(\mem<4><8> ), .B(n148), .Y(n1711) );
  OAI21X1 U1678 ( .A(n147), .B(n1233), .C(n1711), .Y(n1859) );
  NAND2X1 U1679 ( .A(\mem<4><9> ), .B(n148), .Y(n1712) );
  OAI21X1 U1680 ( .A(n147), .B(n1235), .C(n1712), .Y(n1858) );
  NAND2X1 U1681 ( .A(\mem<4><10> ), .B(n148), .Y(n1713) );
  OAI21X1 U1682 ( .A(n147), .B(n1237), .C(n1713), .Y(n1857) );
  NAND2X1 U1683 ( .A(\mem<4><11> ), .B(n148), .Y(n1714) );
  OAI21X1 U1684 ( .A(n147), .B(n1239), .C(n1714), .Y(n1856) );
  NAND2X1 U1685 ( .A(\mem<4><12> ), .B(n148), .Y(n1715) );
  OAI21X1 U1686 ( .A(n147), .B(n1241), .C(n1715), .Y(n1855) );
  NAND2X1 U1687 ( .A(\mem<4><13> ), .B(n148), .Y(n1716) );
  OAI21X1 U1688 ( .A(n147), .B(n1243), .C(n1716), .Y(n1854) );
  NAND2X1 U1689 ( .A(\mem<4><14> ), .B(n148), .Y(n1717) );
  OAI21X1 U1690 ( .A(n147), .B(n1245), .C(n1717), .Y(n1853) );
  NAND2X1 U1691 ( .A(\mem<4><15> ), .B(n148), .Y(n1718) );
  OAI21X1 U1692 ( .A(n147), .B(n1247), .C(n1718), .Y(n1852) );
  NAND2X1 U1693 ( .A(\mem<3><0> ), .B(n151), .Y(n1720) );
  OAI21X1 U1694 ( .A(n150), .B(n1217), .C(n1720), .Y(n1851) );
  NAND2X1 U1695 ( .A(\mem<3><1> ), .B(n151), .Y(n1721) );
  OAI21X1 U1696 ( .A(n150), .B(n1219), .C(n1721), .Y(n1850) );
  NAND2X1 U1697 ( .A(\mem<3><2> ), .B(n151), .Y(n1722) );
  OAI21X1 U1698 ( .A(n150), .B(n1221), .C(n1722), .Y(n1849) );
  NAND2X1 U1699 ( .A(\mem<3><3> ), .B(n151), .Y(n1723) );
  OAI21X1 U1700 ( .A(n150), .B(n1223), .C(n1723), .Y(n1848) );
  NAND2X1 U1701 ( .A(\mem<3><4> ), .B(n151), .Y(n1724) );
  OAI21X1 U1702 ( .A(n150), .B(n1225), .C(n1724), .Y(n1847) );
  NAND2X1 U1703 ( .A(\mem<3><5> ), .B(n151), .Y(n1725) );
  OAI21X1 U1704 ( .A(n150), .B(n1227), .C(n1725), .Y(n1846) );
  NAND2X1 U1705 ( .A(\mem<3><6> ), .B(n151), .Y(n1726) );
  OAI21X1 U1706 ( .A(n150), .B(n1229), .C(n1726), .Y(n1845) );
  NAND2X1 U1707 ( .A(\mem<3><7> ), .B(n151), .Y(n1727) );
  OAI21X1 U1708 ( .A(n150), .B(n1231), .C(n1727), .Y(n1844) );
  NAND2X1 U1709 ( .A(\mem<3><8> ), .B(n151), .Y(n1728) );
  OAI21X1 U1710 ( .A(n150), .B(n1233), .C(n1728), .Y(n1843) );
  NAND2X1 U1711 ( .A(\mem<3><9> ), .B(n151), .Y(n1729) );
  OAI21X1 U1712 ( .A(n150), .B(n1235), .C(n1729), .Y(n1842) );
  NAND2X1 U1713 ( .A(\mem<3><10> ), .B(n151), .Y(n1730) );
  OAI21X1 U1714 ( .A(n150), .B(n1237), .C(n1730), .Y(n1841) );
  NAND2X1 U1715 ( .A(\mem<3><11> ), .B(n151), .Y(n1731) );
  OAI21X1 U1716 ( .A(n150), .B(n1239), .C(n1731), .Y(n1840) );
  NAND2X1 U1717 ( .A(\mem<3><12> ), .B(n151), .Y(n1732) );
  OAI21X1 U1718 ( .A(n150), .B(n1241), .C(n1732), .Y(n1839) );
  NAND2X1 U1719 ( .A(\mem<3><13> ), .B(n151), .Y(n1733) );
  OAI21X1 U1720 ( .A(n150), .B(n1243), .C(n1733), .Y(n1838) );
  NAND2X1 U1721 ( .A(\mem<3><14> ), .B(n151), .Y(n1734) );
  OAI21X1 U1722 ( .A(n150), .B(n1245), .C(n1734), .Y(n1837) );
  NAND2X1 U1723 ( .A(\mem<3><15> ), .B(n151), .Y(n1735) );
  OAI21X1 U1724 ( .A(n150), .B(n1247), .C(n1735), .Y(n1836) );
  NAND2X1 U1725 ( .A(\mem<2><0> ), .B(n154), .Y(n1737) );
  OAI21X1 U1726 ( .A(n153), .B(n1218), .C(n1737), .Y(n1835) );
  NAND2X1 U1727 ( .A(\mem<2><1> ), .B(n154), .Y(n1738) );
  OAI21X1 U1728 ( .A(n153), .B(n1219), .C(n1738), .Y(n1834) );
  NAND2X1 U1729 ( .A(\mem<2><2> ), .B(n154), .Y(n1739) );
  OAI21X1 U1730 ( .A(n153), .B(n1221), .C(n1739), .Y(n1833) );
  NAND2X1 U1731 ( .A(\mem<2><3> ), .B(n154), .Y(n1740) );
  OAI21X1 U1732 ( .A(n153), .B(n1223), .C(n1740), .Y(n1832) );
  NAND2X1 U1733 ( .A(\mem<2><4> ), .B(n154), .Y(n1741) );
  OAI21X1 U1734 ( .A(n153), .B(n1225), .C(n1741), .Y(n1831) );
  NAND2X1 U1735 ( .A(\mem<2><5> ), .B(n154), .Y(n1742) );
  OAI21X1 U1736 ( .A(n153), .B(n1227), .C(n1742), .Y(n1830) );
  NAND2X1 U1737 ( .A(\mem<2><6> ), .B(n154), .Y(n1743) );
  OAI21X1 U1738 ( .A(n153), .B(n1229), .C(n1743), .Y(n1829) );
  NAND2X1 U1739 ( .A(\mem<2><7> ), .B(n154), .Y(n1744) );
  OAI21X1 U1740 ( .A(n153), .B(n1231), .C(n1744), .Y(n1828) );
  NAND2X1 U1741 ( .A(\mem<2><8> ), .B(n154), .Y(n1745) );
  OAI21X1 U1742 ( .A(n153), .B(n1233), .C(n1745), .Y(n1827) );
  NAND2X1 U1743 ( .A(\mem<2><9> ), .B(n154), .Y(n1746) );
  OAI21X1 U1744 ( .A(n153), .B(n1235), .C(n1746), .Y(n1826) );
  NAND2X1 U1745 ( .A(\mem<2><10> ), .B(n154), .Y(n1747) );
  OAI21X1 U1746 ( .A(n153), .B(n1237), .C(n1747), .Y(n1825) );
  NAND2X1 U1747 ( .A(\mem<2><11> ), .B(n154), .Y(n1748) );
  OAI21X1 U1748 ( .A(n153), .B(n1239), .C(n1748), .Y(n1824) );
  NAND2X1 U1749 ( .A(\mem<2><12> ), .B(n154), .Y(n1749) );
  OAI21X1 U1750 ( .A(n153), .B(n1241), .C(n1749), .Y(n1823) );
  NAND2X1 U1751 ( .A(\mem<2><13> ), .B(n154), .Y(n1750) );
  OAI21X1 U1752 ( .A(n153), .B(n1243), .C(n1750), .Y(n1822) );
  NAND2X1 U1753 ( .A(\mem<2><14> ), .B(n154), .Y(n1751) );
  OAI21X1 U1754 ( .A(n153), .B(n1245), .C(n1751), .Y(n1821) );
  NAND2X1 U1755 ( .A(\mem<2><15> ), .B(n154), .Y(n1752) );
  OAI21X1 U1756 ( .A(n153), .B(n1247), .C(n1752), .Y(n1820) );
  NAND2X1 U1757 ( .A(\mem<1><0> ), .B(n157), .Y(n1754) );
  OAI21X1 U1758 ( .A(n156), .B(n1217), .C(n1754), .Y(n1819) );
  NAND2X1 U1759 ( .A(\mem<1><1> ), .B(n157), .Y(n1755) );
  OAI21X1 U1760 ( .A(n156), .B(n1219), .C(n1755), .Y(n1818) );
  NAND2X1 U1761 ( .A(\mem<1><2> ), .B(n157), .Y(n1756) );
  OAI21X1 U1762 ( .A(n156), .B(n1221), .C(n1756), .Y(n1817) );
  NAND2X1 U1763 ( .A(\mem<1><3> ), .B(n157), .Y(n1757) );
  OAI21X1 U1764 ( .A(n156), .B(n1223), .C(n1757), .Y(n1816) );
  NAND2X1 U1765 ( .A(\mem<1><4> ), .B(n157), .Y(n1758) );
  OAI21X1 U1766 ( .A(n156), .B(n1225), .C(n1758), .Y(n1815) );
  NAND2X1 U1767 ( .A(\mem<1><5> ), .B(n157), .Y(n1759) );
  OAI21X1 U1768 ( .A(n156), .B(n1227), .C(n1759), .Y(n1814) );
  NAND2X1 U1769 ( .A(\mem<1><6> ), .B(n157), .Y(n1760) );
  OAI21X1 U1770 ( .A(n156), .B(n1229), .C(n1760), .Y(n1813) );
  NAND2X1 U1771 ( .A(\mem<1><7> ), .B(n157), .Y(n1761) );
  OAI21X1 U1772 ( .A(n156), .B(n1231), .C(n1761), .Y(n1812) );
  NAND2X1 U1773 ( .A(\mem<1><8> ), .B(n157), .Y(n1762) );
  OAI21X1 U1774 ( .A(n156), .B(n1233), .C(n1762), .Y(n1811) );
  NAND2X1 U1775 ( .A(\mem<1><9> ), .B(n157), .Y(n1763) );
  OAI21X1 U1776 ( .A(n156), .B(n1235), .C(n1763), .Y(n1810) );
  NAND2X1 U1777 ( .A(\mem<1><10> ), .B(n157), .Y(n1764) );
  OAI21X1 U1778 ( .A(n156), .B(n1237), .C(n1764), .Y(n1809) );
  NAND2X1 U1779 ( .A(\mem<1><11> ), .B(n157), .Y(n1765) );
  OAI21X1 U1780 ( .A(n156), .B(n1239), .C(n1765), .Y(n1808) );
  NAND2X1 U1781 ( .A(\mem<1><12> ), .B(n157), .Y(n1766) );
  OAI21X1 U1782 ( .A(n156), .B(n1241), .C(n1766), .Y(n1807) );
  NAND2X1 U1783 ( .A(\mem<1><13> ), .B(n157), .Y(n1767) );
  OAI21X1 U1784 ( .A(n156), .B(n1243), .C(n1767), .Y(n1806) );
  NAND2X1 U1785 ( .A(\mem<1><14> ), .B(n157), .Y(n1768) );
  OAI21X1 U1786 ( .A(n156), .B(n1245), .C(n1768), .Y(n1805) );
  NAND2X1 U1787 ( .A(\mem<1><15> ), .B(n157), .Y(n1769) );
  OAI21X1 U1788 ( .A(n156), .B(n1247), .C(n1769), .Y(n1804) );
  NAND2X1 U1789 ( .A(\mem<0><0> ), .B(n158), .Y(n1772) );
  OAI21X1 U1790 ( .A(n70), .B(n1218), .C(n1772), .Y(n1803) );
  NAND2X1 U1791 ( .A(\mem<0><1> ), .B(n158), .Y(n1773) );
  OAI21X1 U1792 ( .A(n70), .B(n1219), .C(n1773), .Y(n1802) );
  NAND2X1 U1793 ( .A(\mem<0><2> ), .B(n158), .Y(n1774) );
  OAI21X1 U1794 ( .A(n70), .B(n1221), .C(n1774), .Y(n1801) );
  NAND2X1 U1795 ( .A(\mem<0><3> ), .B(n158), .Y(n1775) );
  OAI21X1 U1796 ( .A(n70), .B(n1223), .C(n1775), .Y(n1800) );
  NAND2X1 U1797 ( .A(\mem<0><4> ), .B(n158), .Y(n1776) );
  OAI21X1 U1798 ( .A(n70), .B(n1225), .C(n1776), .Y(n1799) );
  NAND2X1 U1799 ( .A(\mem<0><5> ), .B(n158), .Y(n1777) );
  OAI21X1 U1800 ( .A(n70), .B(n1227), .C(n1777), .Y(n1798) );
  NAND2X1 U1801 ( .A(\mem<0><6> ), .B(n158), .Y(n1778) );
  OAI21X1 U1802 ( .A(n70), .B(n1229), .C(n1778), .Y(n1797) );
  NAND2X1 U1803 ( .A(\mem<0><7> ), .B(n158), .Y(n1779) );
  OAI21X1 U1804 ( .A(n70), .B(n1231), .C(n1779), .Y(n1796) );
  NAND2X1 U1805 ( .A(\mem<0><8> ), .B(n158), .Y(n1780) );
  OAI21X1 U1806 ( .A(n70), .B(n1233), .C(n1780), .Y(n1795) );
  NAND2X1 U1807 ( .A(\mem<0><9> ), .B(n158), .Y(n1781) );
  OAI21X1 U1808 ( .A(n70), .B(n1235), .C(n1781), .Y(n1794) );
  NAND2X1 U1809 ( .A(\mem<0><10> ), .B(n158), .Y(n1782) );
  OAI21X1 U1810 ( .A(n70), .B(n1237), .C(n1782), .Y(n1793) );
  NAND2X1 U1811 ( .A(\mem<0><11> ), .B(n158), .Y(n1783) );
  OAI21X1 U1812 ( .A(n70), .B(n1239), .C(n1783), .Y(n1792) );
  NAND2X1 U1813 ( .A(\mem<0><12> ), .B(n158), .Y(n1784) );
  OAI21X1 U1814 ( .A(n70), .B(n1241), .C(n1784), .Y(n1791) );
  NAND2X1 U1815 ( .A(\mem<0><13> ), .B(n158), .Y(n1785) );
  OAI21X1 U1816 ( .A(n70), .B(n1243), .C(n1785), .Y(n1790) );
  NAND2X1 U1817 ( .A(\mem<0><14> ), .B(n158), .Y(n1786) );
  OAI21X1 U1818 ( .A(n70), .B(n1245), .C(n1786), .Y(n1789) );
  NAND2X1 U1819 ( .A(\mem<0><15> ), .B(n158), .Y(n1787) );
  OAI21X1 U1820 ( .A(n70), .B(n1247), .C(n1787), .Y(n1788) );
endmodule


module memc_Size16_0 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n1832), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n1833), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n1834), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n1835), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n1836), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n1837), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n1838), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n1839), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n1840), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1841), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1842), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1843), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1844), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1845), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1846), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1847), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n1848), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n1849), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n1850), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n1851), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n1852), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n1853), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n1854), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n1855), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1856), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1857), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1858), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1859), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1860), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1861), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1862), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1863), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n1864), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n1865), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n1866), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n1867), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n1868), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n1869), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n1870), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n1871), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1872), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1873), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1874), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1875), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1876), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1877), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1878), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1879), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n1880), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n1881), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n1882), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n1883), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n1884), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n1885), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n1886), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n1887), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1888), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1889), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1890), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1891), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1892), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1893), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1894), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1895), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n1896), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n1897), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n1898), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n1899), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n1900), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n1901), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n1902), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n1903), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1904), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1905), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1906), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1907), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1908), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1909), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1910), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1911), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n1912), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n1913), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n1914), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n1915), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n1916), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n1917), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n1918), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n1919), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1920), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1921), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1922), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1923), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1924), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1925), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1926), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1927), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n1928), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n1929), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n1930), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n1931), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n1932), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n1933), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n1934), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n1935), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1936), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1937), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1938), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1939), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1940), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1941), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1942), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1943), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n1944), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n1945), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n1946), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n1947), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n1948), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n1949), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n1950), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n1951), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1952), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1953), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1954), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1955), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1956), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1957), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1958), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1959), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n1960), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n1961), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n1962), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n1963), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n1964), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n1965), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n1966), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n1967), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1968), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1969), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1970), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1971), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1972), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1973), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1974), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1975), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n1976), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n1977), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n1978), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n1979), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n1980), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n1981), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n1982), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n1983), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n1984), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n1985), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n1986), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n1987), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n1988), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n1989), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n1990), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n1991), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n1992), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n1993), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n1994), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n1995), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n1996), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n1997), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n1998), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n1999), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n2000), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n2001), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n2002), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n2003), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n2004), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n2005), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n2006), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n2007), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n2008), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n2009), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n2010), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n2011), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n2012), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n2013), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n2014), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n2015), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n2016), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n2017), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n2018), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n2019), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n2020), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n2021), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n2022), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n2023), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n2024), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n2025), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n2026), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n2027), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n2028), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n2029), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n2030), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n2031), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2032), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2033), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2034), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2035), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2036), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2037), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2038), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2039), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n2040), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n2041), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n2042), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n2043), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n2044), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n2045), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n2046), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n2047), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2048), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2049), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2050), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2051), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2052), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2053), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2054), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2055), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n2056), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n2057), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n2058), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n2059), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n2060), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n2061), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n2062), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n2063), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2064), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2065), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2066), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2067), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2068), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2069), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2070), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2071), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n2072), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n2073), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n2074), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n2075), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n2076), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n2077), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n2078), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n2079), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2080), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2081), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2082), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2083), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2084), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2085), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2086), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2087), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n2088), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n2089), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n2090), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n2091), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n2092), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n2093), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n2094), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n2095), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2096), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2097), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2098), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2099), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2100), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2101), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2102), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2103), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n2104), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n2105), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n2106), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n2107), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n2108), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n2109), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n2110), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n2111), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2112), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2113), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2114), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2115), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2116), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2117), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2118), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2119), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n2120), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n2121), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n2122), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n2123), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n2124), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n2125), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n2126), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n2127), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2128), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2129), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2130), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2131), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2132), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2133), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2134), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2135), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n2136), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n2137), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n2138), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n2139), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n2140), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n2141), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n2142), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n2143), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2144), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2145), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2146), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2147), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2148), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2149), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2150), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2151), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n2152), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n2153), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n2154), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n2155), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n2156), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n2157), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n2158), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n2159), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2160), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2161), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2162), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2163), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2164), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2165), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2166), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2167), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n2168), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n2169), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n2170), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n2171), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n2172), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n2173), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n2174), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n2175), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2176), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2177), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2178), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2179), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2180), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2181), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2182), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2183), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n2184), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n2185), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n2186), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n2187), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n2188), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n2189), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n2190), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n2191), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2192), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2193), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2194), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2195), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2196), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2197), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2198), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2199), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n2200), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n2201), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n2202), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n2203), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n2204), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n2205), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n2206), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n2207), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2208), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2209), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2210), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2211), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2212), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2213), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2214), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2215), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n2216), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n2217), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n2218), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n2219), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n2220), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n2221), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n2222), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n2223), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2224), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2225), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2226), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2227), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2228), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2229), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2230), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2231), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n2232), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n2233), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n2234), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n2235), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n2236), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n2237), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n2238), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n2239), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2240), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2241), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2242), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2243), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2244), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2245), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2246), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2247), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n2248), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n2249), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n2250), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n2251), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n2252), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n2253), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n2254), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n2255), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2256), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2257), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2258), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2259), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2260), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2261), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2262), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2263), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n2264), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n2265), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n2266), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n2267), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n2268), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n2269), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n2270), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n2271), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2272), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2273), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2274), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2275), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2276), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2277), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2278), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2279), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n2280), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n2281), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n2282), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n2283), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n2284), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n2285), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n2286), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n2287), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2288), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2289), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2290), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2291), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2292), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2293), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2294), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2295), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n2296), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n2297), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n2298), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n2299), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n2300), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n2301), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n2302), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n2303), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2304), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2305), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2306), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2307), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2308), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2309), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2310), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2311), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n2312), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n2313), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n2314), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n2315), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n2316), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n2317), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n2318), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n2319), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2320), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2321), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2322), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2323), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2324), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2325), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2326), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2327), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n2328), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n2329), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n2330), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n2331), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n2332), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n2333), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n2334), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n2335), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2336), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2337), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2338), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2339), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2340), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2341), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2342), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2343), .CLK(clk), .Q(\mem<31><0> ) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n2344) );
  INVX2 U2 ( .A(N10), .Y(n1296) );
  INVX1 U3 ( .A(n1296), .Y(n1205) );
  INVX1 U4 ( .A(n1194), .Y(n1203) );
  INVX1 U5 ( .A(n1194), .Y(n1204) );
  INVX1 U6 ( .A(n1194), .Y(n1211) );
  INVX1 U7 ( .A(n1195), .Y(n1210) );
  INVX1 U8 ( .A(n1212), .Y(n1195) );
  INVX1 U9 ( .A(n1296), .Y(n1196) );
  INVX4 U10 ( .A(n54), .Y(n143) );
  INVX4 U11 ( .A(n53), .Y(n140) );
  INVX1 U12 ( .A(n1166), .Y(N23) );
  INVX1 U13 ( .A(n1169), .Y(N20) );
  INVX1 U14 ( .A(n1212), .Y(n1194) );
  INVX1 U15 ( .A(n1193), .Y(n1182) );
  INVX1 U16 ( .A(n1193), .Y(n1183) );
  INVX2 U17 ( .A(n1195), .Y(n1197) );
  INVX1 U18 ( .A(n1193), .Y(n1184) );
  INVX2 U19 ( .A(n1195), .Y(n1198) );
  INVX1 U20 ( .A(n1181), .Y(n1185) );
  INVX2 U21 ( .A(n1195), .Y(n1200) );
  INVX1 U22 ( .A(n1181), .Y(n1186) );
  INVX2 U23 ( .A(n1195), .Y(n1201) );
  INVX1 U24 ( .A(n1181), .Y(n1187) );
  INVX1 U25 ( .A(n1180), .Y(n1188) );
  INVX2 U26 ( .A(n1194), .Y(n1206) );
  INVX1 U27 ( .A(n1180), .Y(n1189) );
  INVX2 U28 ( .A(n1194), .Y(n1207) );
  INVX2 U29 ( .A(n1194), .Y(n1208) );
  INVX1 U30 ( .A(n1180), .Y(n1190) );
  INVX2 U31 ( .A(n1195), .Y(n1209) );
  INVX1 U32 ( .A(n1181), .Y(n1191) );
  INVX2 U33 ( .A(n1194), .Y(n1199) );
  INVX1 U34 ( .A(n1180), .Y(n1192) );
  INVX1 U35 ( .A(n645), .Y(N32) );
  INVX1 U36 ( .A(n646), .Y(N31) );
  INVX1 U37 ( .A(n647), .Y(N30) );
  INVX1 U38 ( .A(n648), .Y(N29) );
  INVX1 U39 ( .A(n649), .Y(N28) );
  INVX1 U40 ( .A(n650), .Y(N27) );
  INVX1 U41 ( .A(n1163), .Y(N26) );
  INVX1 U42 ( .A(n1164), .Y(N25) );
  INVX1 U43 ( .A(n1165), .Y(N24) );
  INVX1 U44 ( .A(n1167), .Y(N22) );
  INVX1 U45 ( .A(n1168), .Y(N21) );
  INVX1 U46 ( .A(n1170), .Y(N19) );
  INVX1 U47 ( .A(n1171), .Y(N18) );
  INVX1 U48 ( .A(n1172), .Y(N17) );
  INVX1 U49 ( .A(n1299), .Y(n1178) );
  INVX1 U50 ( .A(n1299), .Y(n1179) );
  INVX2 U51 ( .A(n1195), .Y(n1202) );
  INVX1 U52 ( .A(N14), .Y(n1302) );
  INVX1 U53 ( .A(n1297), .Y(n1193) );
  INVX1 U54 ( .A(n1299), .Y(n1177) );
  INVX1 U55 ( .A(n1299), .Y(n1176) );
  INVX1 U56 ( .A(n1300), .Y(n1174) );
  INVX1 U57 ( .A(n1300), .Y(n1175) );
  INVX1 U58 ( .A(n1297), .Y(n1181) );
  INVX1 U59 ( .A(n1297), .Y(n1180) );
  INVX1 U60 ( .A(n1302), .Y(n1173) );
  INVX1 U61 ( .A(rst), .Y(n1295) );
  INVX1 U62 ( .A(n92), .Y(n1227) );
  INVX1 U63 ( .A(n93), .Y(n1244) );
  INVX1 U64 ( .A(n94), .Y(n1261) );
  INVX1 U65 ( .A(n95), .Y(n1264) );
  INVX4 U66 ( .A(n62), .Y(n1270) );
  INVX1 U67 ( .A(write), .Y(n1) );
  INVX1 U68 ( .A(n1), .Y(n2) );
  INVX1 U69 ( .A(n1303), .Y(n1304) );
  INVX2 U70 ( .A(n1303), .Y(n4) );
  INVX1 U71 ( .A(n1303), .Y(n3) );
  INVX1 U72 ( .A(N13), .Y(n1300) );
  AND2X2 U73 ( .A(n1267), .B(n96), .Y(n5) );
  INVX1 U74 ( .A(n5), .Y(n6) );
  AND2X2 U75 ( .A(n1269), .B(n98), .Y(n7) );
  INVX1 U76 ( .A(n7), .Y(n8) );
  AND2X2 U77 ( .A(n1267), .B(n100), .Y(n9) );
  INVX1 U78 ( .A(n9), .Y(n10) );
  AND2X2 U79 ( .A(n1269), .B(n102), .Y(n11) );
  INVX1 U80 ( .A(n11), .Y(n12) );
  AND2X2 U81 ( .A(n1267), .B(n104), .Y(n13) );
  INVX1 U82 ( .A(n13), .Y(n14) );
  AND2X2 U83 ( .A(n1269), .B(n106), .Y(n15) );
  INVX1 U84 ( .A(n15), .Y(n16) );
  AND2X2 U85 ( .A(n1268), .B(n108), .Y(n17) );
  INVX1 U86 ( .A(n17), .Y(n18) );
  AND2X2 U87 ( .A(n1269), .B(n92), .Y(n19) );
  INVX1 U88 ( .A(n19), .Y(n20) );
  AND2X2 U89 ( .A(n1267), .B(n110), .Y(n21) );
  INVX1 U90 ( .A(n21), .Y(n22) );
  AND2X2 U91 ( .A(n1269), .B(n112), .Y(n23) );
  INVX1 U92 ( .A(n23), .Y(n24) );
  AND2X2 U93 ( .A(n1268), .B(n114), .Y(n25) );
  INVX1 U94 ( .A(n25), .Y(n26) );
  AND2X2 U95 ( .A(n1267), .B(n116), .Y(n27) );
  INVX1 U96 ( .A(n27), .Y(n28) );
  AND2X2 U97 ( .A(n1267), .B(n118), .Y(n29) );
  INVX1 U98 ( .A(n29), .Y(n30) );
  AND2X2 U99 ( .A(n1267), .B(n120), .Y(n31) );
  INVX1 U100 ( .A(n31), .Y(n32) );
  AND2X2 U101 ( .A(n1267), .B(n122), .Y(n33) );
  INVX1 U102 ( .A(n33), .Y(n34) );
  AND2X2 U103 ( .A(n1267), .B(n93), .Y(n35) );
  INVX1 U104 ( .A(n35), .Y(n36) );
  AND2X2 U105 ( .A(n1267), .B(n124), .Y(n37) );
  INVX1 U106 ( .A(n37), .Y(n38) );
  AND2X2 U107 ( .A(n1267), .B(n126), .Y(n39) );
  INVX1 U108 ( .A(n39), .Y(n40) );
  AND2X2 U109 ( .A(n1267), .B(n128), .Y(n41) );
  INVX1 U110 ( .A(n41), .Y(n42) );
  AND2X2 U111 ( .A(n1267), .B(n130), .Y(n43) );
  INVX1 U112 ( .A(n43), .Y(n44) );
  AND2X2 U113 ( .A(n1267), .B(n132), .Y(n45) );
  INVX1 U114 ( .A(n45), .Y(n46) );
  AND2X2 U115 ( .A(n1267), .B(n134), .Y(n47) );
  INVX1 U116 ( .A(n47), .Y(n48) );
  AND2X2 U117 ( .A(n1267), .B(n136), .Y(n49) );
  INVX1 U118 ( .A(n49), .Y(n50) );
  AND2X2 U119 ( .A(n1268), .B(n94), .Y(n51) );
  INVX1 U120 ( .A(n51), .Y(n52) );
  AND2X2 U121 ( .A(n1268), .B(n138), .Y(n53) );
  AND2X2 U122 ( .A(n1268), .B(n141), .Y(n54) );
  AND2X2 U123 ( .A(n1268), .B(n144), .Y(n55) );
  AND2X2 U124 ( .A(n1268), .B(n148), .Y(n56) );
  AND2X2 U125 ( .A(n1268), .B(n152), .Y(n57) );
  AND2X2 U126 ( .A(n1268), .B(n156), .Y(n58) );
  AND2X2 U127 ( .A(n1268), .B(n160), .Y(n59) );
  AND2X2 U128 ( .A(n1267), .B(n95), .Y(n60) );
  INVX1 U129 ( .A(n60), .Y(n61) );
  BUFX2 U130 ( .A(n6), .Y(n1213) );
  BUFX2 U131 ( .A(n6), .Y(n1214) );
  BUFX2 U132 ( .A(n8), .Y(n1215) );
  BUFX2 U133 ( .A(n8), .Y(n1216) );
  BUFX2 U134 ( .A(n10), .Y(n1217) );
  BUFX2 U135 ( .A(n10), .Y(n1218) );
  BUFX2 U136 ( .A(n12), .Y(n1219) );
  BUFX2 U137 ( .A(n12), .Y(n1220) );
  BUFX2 U138 ( .A(n14), .Y(n1221) );
  BUFX2 U139 ( .A(n14), .Y(n1222) );
  BUFX2 U140 ( .A(n16), .Y(n1223) );
  BUFX2 U141 ( .A(n16), .Y(n1224) );
  BUFX2 U142 ( .A(n18), .Y(n1225) );
  BUFX2 U143 ( .A(n18), .Y(n1226) );
  BUFX2 U144 ( .A(n20), .Y(n1228) );
  BUFX2 U145 ( .A(n20), .Y(n1229) );
  BUFX2 U146 ( .A(n22), .Y(n1230) );
  BUFX2 U147 ( .A(n22), .Y(n1231) );
  BUFX2 U148 ( .A(n24), .Y(n1232) );
  BUFX2 U149 ( .A(n24), .Y(n1233) );
  BUFX2 U150 ( .A(n26), .Y(n1234) );
  BUFX2 U151 ( .A(n26), .Y(n1235) );
  BUFX2 U152 ( .A(n28), .Y(n1236) );
  BUFX2 U153 ( .A(n28), .Y(n1237) );
  BUFX2 U154 ( .A(n30), .Y(n1238) );
  BUFX2 U155 ( .A(n30), .Y(n1239) );
  BUFX2 U156 ( .A(n32), .Y(n1240) );
  BUFX2 U157 ( .A(n32), .Y(n1241) );
  BUFX2 U158 ( .A(n34), .Y(n1242) );
  BUFX2 U159 ( .A(n34), .Y(n1243) );
  BUFX2 U160 ( .A(n36), .Y(n1245) );
  BUFX2 U161 ( .A(n36), .Y(n1246) );
  BUFX2 U162 ( .A(n38), .Y(n1247) );
  BUFX2 U163 ( .A(n38), .Y(n1248) );
  BUFX2 U164 ( .A(n40), .Y(n1249) );
  BUFX2 U165 ( .A(n40), .Y(n1250) );
  BUFX2 U166 ( .A(n42), .Y(n1251) );
  BUFX2 U167 ( .A(n42), .Y(n1252) );
  BUFX2 U168 ( .A(n44), .Y(n1253) );
  BUFX2 U169 ( .A(n44), .Y(n1254) );
  BUFX2 U170 ( .A(n46), .Y(n1255) );
  BUFX2 U171 ( .A(n46), .Y(n1256) );
  BUFX2 U172 ( .A(n48), .Y(n1257) );
  BUFX2 U173 ( .A(n48), .Y(n1258) );
  BUFX2 U174 ( .A(n50), .Y(n1259) );
  BUFX2 U175 ( .A(n50), .Y(n1260) );
  BUFX2 U176 ( .A(n52), .Y(n1262) );
  BUFX2 U177 ( .A(n52), .Y(n1263) );
  BUFX2 U178 ( .A(n61), .Y(n1265) );
  BUFX2 U179 ( .A(n61), .Y(n1266) );
  AND2X2 U180 ( .A(n2), .B(n1295), .Y(n62) );
  INVX1 U181 ( .A(n1298), .Y(n1297) );
  AND2X1 U182 ( .A(n1177), .B(n1297), .Y(n63) );
  AND2X1 U183 ( .A(n2344), .B(n1301), .Y(n64) );
  INVX1 U184 ( .A(n1302), .Y(n1301) );
  BUFX2 U185 ( .A(n1337), .Y(n65) );
  INVX1 U186 ( .A(n65), .Y(n1729) );
  BUFX2 U187 ( .A(n1354), .Y(n66) );
  INVX1 U188 ( .A(n66), .Y(n1746) );
  BUFX2 U189 ( .A(n1371), .Y(n67) );
  INVX1 U190 ( .A(n67), .Y(n1763) );
  BUFX2 U191 ( .A(n1388), .Y(n68) );
  INVX1 U192 ( .A(n68), .Y(n1780) );
  BUFX2 U193 ( .A(n1405), .Y(n69) );
  INVX1 U194 ( .A(n69), .Y(n1797) );
  BUFX2 U195 ( .A(n1566), .Y(n70) );
  INVX1 U196 ( .A(n70), .Y(n1679) );
  BUFX2 U197 ( .A(n1696), .Y(n71) );
  INVX1 U198 ( .A(n71), .Y(n1814) );
  AND2X1 U199 ( .A(n1196), .B(n63), .Y(n72) );
  AND2X1 U200 ( .A(n1175), .B(n64), .Y(n73) );
  AND2X1 U201 ( .A(n1296), .B(n63), .Y(n74) );
  AND2X1 U202 ( .A(n1300), .B(n64), .Y(n75) );
  AND2X2 U203 ( .A(\data_in<0> ), .B(n1269), .Y(n76) );
  AND2X2 U204 ( .A(\data_in<1> ), .B(n1269), .Y(n77) );
  AND2X2 U205 ( .A(\data_in<2> ), .B(n1269), .Y(n78) );
  AND2X2 U206 ( .A(\data_in<3> ), .B(n1269), .Y(n79) );
  AND2X2 U207 ( .A(\data_in<4> ), .B(n1269), .Y(n80) );
  AND2X2 U208 ( .A(\data_in<5> ), .B(n1269), .Y(n81) );
  AND2X2 U209 ( .A(\data_in<6> ), .B(n1269), .Y(n82) );
  AND2X2 U210 ( .A(\data_in<7> ), .B(n1269), .Y(n83) );
  AND2X2 U211 ( .A(\data_in<8> ), .B(n1269), .Y(n84) );
  AND2X2 U212 ( .A(\data_in<9> ), .B(n1269), .Y(n85) );
  AND2X2 U213 ( .A(\data_in<10> ), .B(n1269), .Y(n86) );
  AND2X2 U214 ( .A(\data_in<11> ), .B(n1268), .Y(n87) );
  AND2X2 U215 ( .A(\data_in<12> ), .B(n1268), .Y(n88) );
  AND2X2 U216 ( .A(\data_in<13> ), .B(n1268), .Y(n89) );
  AND2X2 U217 ( .A(\data_in<14> ), .B(n1268), .Y(n90) );
  AND2X2 U218 ( .A(\data_in<15> ), .B(n1268), .Y(n91) );
  AND2X1 U219 ( .A(n73), .B(n1815), .Y(n92) );
  AND2X1 U220 ( .A(n1815), .B(n75), .Y(n93) );
  AND2X1 U221 ( .A(n1815), .B(n1679), .Y(n94) );
  AND2X1 U222 ( .A(n1815), .B(n1814), .Y(n95) );
  AND2X1 U223 ( .A(n72), .B(n73), .Y(n96) );
  INVX1 U224 ( .A(n96), .Y(n97) );
  AND2X1 U225 ( .A(n73), .B(n74), .Y(n98) );
  INVX1 U226 ( .A(n98), .Y(n99) );
  AND2X1 U227 ( .A(n73), .B(n1729), .Y(n100) );
  INVX1 U228 ( .A(n100), .Y(n101) );
  AND2X1 U229 ( .A(n73), .B(n1746), .Y(n102) );
  INVX1 U230 ( .A(n102), .Y(n103) );
  AND2X1 U231 ( .A(n73), .B(n1763), .Y(n104) );
  INVX1 U232 ( .A(n104), .Y(n105) );
  AND2X1 U233 ( .A(n73), .B(n1780), .Y(n106) );
  INVX1 U234 ( .A(n106), .Y(n107) );
  AND2X1 U235 ( .A(n73), .B(n1797), .Y(n108) );
  INVX1 U236 ( .A(n108), .Y(n109) );
  AND2X1 U237 ( .A(n72), .B(n75), .Y(n110) );
  INVX1 U238 ( .A(n110), .Y(n111) );
  AND2X1 U239 ( .A(n74), .B(n75), .Y(n112) );
  INVX1 U240 ( .A(n112), .Y(n113) );
  AND2X1 U241 ( .A(n1729), .B(n75), .Y(n114) );
  INVX1 U242 ( .A(n114), .Y(n115) );
  AND2X1 U243 ( .A(n1746), .B(n75), .Y(n116) );
  INVX1 U244 ( .A(n116), .Y(n117) );
  AND2X1 U245 ( .A(n1763), .B(n75), .Y(n118) );
  INVX1 U246 ( .A(n118), .Y(n119) );
  AND2X1 U247 ( .A(n1780), .B(n75), .Y(n120) );
  INVX1 U248 ( .A(n120), .Y(n121) );
  AND2X1 U249 ( .A(n1797), .B(n75), .Y(n122) );
  INVX1 U250 ( .A(n122), .Y(n123) );
  AND2X1 U251 ( .A(n72), .B(n1679), .Y(n124) );
  INVX1 U252 ( .A(n124), .Y(n125) );
  AND2X1 U253 ( .A(n74), .B(n1679), .Y(n126) );
  INVX1 U254 ( .A(n126), .Y(n127) );
  AND2X1 U255 ( .A(n1729), .B(n1679), .Y(n128) );
  INVX1 U256 ( .A(n128), .Y(n129) );
  AND2X1 U257 ( .A(n1746), .B(n1679), .Y(n130) );
  INVX1 U258 ( .A(n130), .Y(n131) );
  AND2X1 U259 ( .A(n1763), .B(n1679), .Y(n132) );
  INVX1 U260 ( .A(n132), .Y(n133) );
  AND2X1 U261 ( .A(n1780), .B(n1679), .Y(n134) );
  INVX1 U262 ( .A(n134), .Y(n135) );
  AND2X1 U263 ( .A(n1797), .B(n1679), .Y(n136) );
  INVX1 U264 ( .A(n136), .Y(n137) );
  AND2X1 U265 ( .A(n72), .B(n1814), .Y(n138) );
  INVX1 U266 ( .A(n138), .Y(n139) );
  AND2X1 U267 ( .A(n74), .B(n1814), .Y(n141) );
  INVX1 U268 ( .A(n141), .Y(n142) );
  AND2X1 U269 ( .A(n1729), .B(n1814), .Y(n144) );
  INVX1 U270 ( .A(n144), .Y(n145) );
  INVX1 U271 ( .A(n55), .Y(n146) );
  INVX1 U272 ( .A(n55), .Y(n147) );
  AND2X1 U273 ( .A(n1746), .B(n1814), .Y(n148) );
  INVX1 U274 ( .A(n148), .Y(n149) );
  INVX1 U275 ( .A(n56), .Y(n150) );
  INVX1 U276 ( .A(n56), .Y(n151) );
  AND2X1 U277 ( .A(n1763), .B(n1814), .Y(n152) );
  INVX1 U278 ( .A(n152), .Y(n153) );
  INVX1 U279 ( .A(n57), .Y(n154) );
  INVX1 U280 ( .A(n57), .Y(n155) );
  AND2X1 U281 ( .A(n1780), .B(n1814), .Y(n156) );
  INVX1 U282 ( .A(n156), .Y(n157) );
  INVX1 U283 ( .A(n58), .Y(n158) );
  INVX1 U284 ( .A(n58), .Y(n159) );
  AND2X1 U285 ( .A(n1797), .B(n1814), .Y(n160) );
  INVX1 U286 ( .A(n160), .Y(n161) );
  INVX1 U287 ( .A(n59), .Y(n162) );
  INVX1 U288 ( .A(n59), .Y(n163) );
  MUX2X1 U289 ( .B(n165), .A(n166), .S(n1182), .Y(n164) );
  MUX2X1 U290 ( .B(n168), .A(n169), .S(n1182), .Y(n167) );
  MUX2X1 U291 ( .B(n171), .A(n172), .S(n1182), .Y(n170) );
  MUX2X1 U292 ( .B(n174), .A(n175), .S(n1182), .Y(n173) );
  MUX2X1 U293 ( .B(n177), .A(n178), .S(n1175), .Y(n176) );
  MUX2X1 U294 ( .B(n180), .A(n181), .S(n1182), .Y(n179) );
  MUX2X1 U295 ( .B(n183), .A(n184), .S(n1182), .Y(n182) );
  MUX2X1 U296 ( .B(n186), .A(n187), .S(n1182), .Y(n185) );
  MUX2X1 U297 ( .B(n189), .A(n190), .S(n1182), .Y(n188) );
  MUX2X1 U298 ( .B(n192), .A(n193), .S(n1175), .Y(n191) );
  MUX2X1 U299 ( .B(n195), .A(n196), .S(n1183), .Y(n194) );
  MUX2X1 U300 ( .B(n198), .A(n199), .S(n1183), .Y(n197) );
  MUX2X1 U301 ( .B(n201), .A(n202), .S(n1183), .Y(n200) );
  MUX2X1 U302 ( .B(n204), .A(n205), .S(n1183), .Y(n203) );
  MUX2X1 U303 ( .B(n207), .A(n208), .S(n1175), .Y(n206) );
  MUX2X1 U304 ( .B(n210), .A(n211), .S(n1183), .Y(n209) );
  MUX2X1 U305 ( .B(n213), .A(n215), .S(n1183), .Y(n212) );
  MUX2X1 U306 ( .B(n217), .A(n218), .S(n1183), .Y(n216) );
  MUX2X1 U307 ( .B(n220), .A(n221), .S(n1183), .Y(n219) );
  MUX2X1 U308 ( .B(n223), .A(n224), .S(n1175), .Y(n222) );
  MUX2X1 U309 ( .B(n226), .A(n227), .S(n1183), .Y(n225) );
  MUX2X1 U310 ( .B(n229), .A(n230), .S(n1183), .Y(n228) );
  MUX2X1 U311 ( .B(n232), .A(n233), .S(n1183), .Y(n231) );
  MUX2X1 U312 ( .B(n235), .A(n236), .S(n1183), .Y(n234) );
  MUX2X1 U313 ( .B(n238), .A(n239), .S(n1175), .Y(n237) );
  MUX2X1 U314 ( .B(n241), .A(n242), .S(n1184), .Y(n240) );
  MUX2X1 U315 ( .B(n244), .A(n245), .S(n1184), .Y(n243) );
  MUX2X1 U316 ( .B(n247), .A(n248), .S(n1184), .Y(n246) );
  MUX2X1 U317 ( .B(n250), .A(n251), .S(n1184), .Y(n249) );
  MUX2X1 U318 ( .B(n253), .A(n254), .S(n1175), .Y(n252) );
  MUX2X1 U319 ( .B(n256), .A(n257), .S(n1184), .Y(n255) );
  MUX2X1 U320 ( .B(n259), .A(n260), .S(n1184), .Y(n258) );
  MUX2X1 U321 ( .B(n262), .A(n263), .S(n1184), .Y(n261) );
  MUX2X1 U322 ( .B(n265), .A(n266), .S(n1184), .Y(n264) );
  MUX2X1 U323 ( .B(n268), .A(n269), .S(n1175), .Y(n267) );
  MUX2X1 U324 ( .B(n271), .A(n272), .S(n1184), .Y(n270) );
  MUX2X1 U325 ( .B(n274), .A(n275), .S(n1184), .Y(n273) );
  MUX2X1 U326 ( .B(n277), .A(n278), .S(n1184), .Y(n276) );
  MUX2X1 U327 ( .B(n280), .A(n281), .S(n1184), .Y(n279) );
  MUX2X1 U328 ( .B(n283), .A(n284), .S(n1175), .Y(n282) );
  MUX2X1 U329 ( .B(n286), .A(n287), .S(n1185), .Y(n285) );
  MUX2X1 U330 ( .B(n289), .A(n290), .S(n1185), .Y(n288) );
  MUX2X1 U331 ( .B(n292), .A(n293), .S(n1185), .Y(n291) );
  MUX2X1 U332 ( .B(n295), .A(n296), .S(n1185), .Y(n294) );
  MUX2X1 U333 ( .B(n298), .A(n299), .S(n1175), .Y(n297) );
  MUX2X1 U334 ( .B(n301), .A(n302), .S(n1185), .Y(n300) );
  MUX2X1 U335 ( .B(n304), .A(n305), .S(n1185), .Y(n303) );
  MUX2X1 U336 ( .B(n307), .A(n308), .S(n1185), .Y(n306) );
  MUX2X1 U337 ( .B(n310), .A(n311), .S(n1185), .Y(n309) );
  MUX2X1 U338 ( .B(n313), .A(n314), .S(n1175), .Y(n312) );
  MUX2X1 U339 ( .B(n316), .A(n317), .S(n1185), .Y(n315) );
  MUX2X1 U340 ( .B(n319), .A(n320), .S(n1185), .Y(n318) );
  MUX2X1 U341 ( .B(n322), .A(n323), .S(n1185), .Y(n321) );
  MUX2X1 U342 ( .B(n325), .A(n326), .S(n1185), .Y(n324) );
  MUX2X1 U343 ( .B(n328), .A(n329), .S(n1175), .Y(n327) );
  MUX2X1 U344 ( .B(n331), .A(n332), .S(n1186), .Y(n330) );
  MUX2X1 U345 ( .B(n334), .A(n335), .S(n1186), .Y(n333) );
  MUX2X1 U346 ( .B(n337), .A(n338), .S(n1186), .Y(n336) );
  MUX2X1 U347 ( .B(n340), .A(n341), .S(n1186), .Y(n339) );
  MUX2X1 U348 ( .B(n343), .A(n344), .S(n1175), .Y(n342) );
  MUX2X1 U349 ( .B(n346), .A(n347), .S(n1186), .Y(n345) );
  MUX2X1 U350 ( .B(n349), .A(n350), .S(n1186), .Y(n348) );
  MUX2X1 U351 ( .B(n352), .A(n353), .S(n1186), .Y(n351) );
  MUX2X1 U352 ( .B(n355), .A(n356), .S(n1186), .Y(n354) );
  MUX2X1 U353 ( .B(n358), .A(n359), .S(n1174), .Y(n357) );
  MUX2X1 U354 ( .B(n361), .A(n362), .S(n1186), .Y(n360) );
  MUX2X1 U355 ( .B(n364), .A(n365), .S(n1186), .Y(n363) );
  MUX2X1 U356 ( .B(n367), .A(n368), .S(n1186), .Y(n366) );
  MUX2X1 U357 ( .B(n370), .A(n371), .S(n1186), .Y(n369) );
  MUX2X1 U358 ( .B(n373), .A(n374), .S(n1174), .Y(n372) );
  MUX2X1 U359 ( .B(n376), .A(n377), .S(n1187), .Y(n375) );
  MUX2X1 U360 ( .B(n379), .A(n380), .S(n1187), .Y(n378) );
  MUX2X1 U361 ( .B(n382), .A(n383), .S(n1187), .Y(n381) );
  MUX2X1 U362 ( .B(n385), .A(n386), .S(n1187), .Y(n384) );
  MUX2X1 U363 ( .B(n388), .A(n389), .S(n1174), .Y(n387) );
  MUX2X1 U364 ( .B(n391), .A(n392), .S(n1187), .Y(n390) );
  MUX2X1 U365 ( .B(n394), .A(n395), .S(n1187), .Y(n393) );
  MUX2X1 U366 ( .B(n397), .A(n398), .S(n1187), .Y(n396) );
  MUX2X1 U367 ( .B(n400), .A(n401), .S(n1187), .Y(n399) );
  MUX2X1 U368 ( .B(n403), .A(n404), .S(n1174), .Y(n402) );
  MUX2X1 U369 ( .B(n406), .A(n407), .S(n1187), .Y(n405) );
  MUX2X1 U370 ( .B(n409), .A(n410), .S(n1187), .Y(n408) );
  MUX2X1 U371 ( .B(n412), .A(n413), .S(n1187), .Y(n411) );
  MUX2X1 U372 ( .B(n415), .A(n416), .S(n1187), .Y(n414) );
  MUX2X1 U373 ( .B(n418), .A(n419), .S(n1174), .Y(n417) );
  MUX2X1 U374 ( .B(n421), .A(n422), .S(n1188), .Y(n420) );
  MUX2X1 U375 ( .B(n424), .A(n425), .S(n1188), .Y(n423) );
  MUX2X1 U376 ( .B(n427), .A(n428), .S(n1188), .Y(n426) );
  MUX2X1 U377 ( .B(n430), .A(n431), .S(n1188), .Y(n429) );
  MUX2X1 U378 ( .B(n433), .A(n434), .S(n1174), .Y(n432) );
  MUX2X1 U379 ( .B(n436), .A(n437), .S(n1188), .Y(n435) );
  MUX2X1 U380 ( .B(n439), .A(n440), .S(n1188), .Y(n438) );
  MUX2X1 U381 ( .B(n442), .A(n443), .S(n1188), .Y(n441) );
  MUX2X1 U382 ( .B(n445), .A(n446), .S(n1188), .Y(n444) );
  MUX2X1 U383 ( .B(n448), .A(n449), .S(n1174), .Y(n447) );
  MUX2X1 U384 ( .B(n451), .A(n452), .S(n1188), .Y(n450) );
  MUX2X1 U385 ( .B(n454), .A(n455), .S(n1188), .Y(n453) );
  MUX2X1 U386 ( .B(n457), .A(n458), .S(n1188), .Y(n456) );
  MUX2X1 U387 ( .B(n460), .A(n461), .S(n1188), .Y(n459) );
  MUX2X1 U388 ( .B(n463), .A(n464), .S(n1174), .Y(n462) );
  MUX2X1 U389 ( .B(n466), .A(n467), .S(n1189), .Y(n465) );
  MUX2X1 U390 ( .B(n469), .A(n470), .S(n1189), .Y(n468) );
  MUX2X1 U391 ( .B(n472), .A(n473), .S(n1189), .Y(n471) );
  MUX2X1 U392 ( .B(n475), .A(n476), .S(n1189), .Y(n474) );
  MUX2X1 U393 ( .B(n478), .A(n479), .S(n1174), .Y(n477) );
  MUX2X1 U394 ( .B(n481), .A(n482), .S(n1189), .Y(n480) );
  MUX2X1 U395 ( .B(n484), .A(n485), .S(n1189), .Y(n483) );
  MUX2X1 U396 ( .B(n487), .A(n488), .S(n1189), .Y(n486) );
  MUX2X1 U397 ( .B(n490), .A(n491), .S(n1189), .Y(n489) );
  MUX2X1 U398 ( .B(n493), .A(n494), .S(n1174), .Y(n492) );
  MUX2X1 U399 ( .B(n496), .A(n497), .S(n1189), .Y(n495) );
  MUX2X1 U400 ( .B(n499), .A(n500), .S(n1189), .Y(n498) );
  MUX2X1 U401 ( .B(n502), .A(n503), .S(n1189), .Y(n501) );
  MUX2X1 U402 ( .B(n505), .A(n506), .S(n1189), .Y(n504) );
  MUX2X1 U403 ( .B(n508), .A(n509), .S(n1174), .Y(n507) );
  MUX2X1 U404 ( .B(n511), .A(n512), .S(n1190), .Y(n510) );
  MUX2X1 U405 ( .B(n514), .A(n515), .S(n1190), .Y(n513) );
  MUX2X1 U406 ( .B(n517), .A(n518), .S(n1190), .Y(n516) );
  MUX2X1 U407 ( .B(n520), .A(n521), .S(n1190), .Y(n519) );
  MUX2X1 U408 ( .B(n523), .A(n524), .S(n1174), .Y(n522) );
  MUX2X1 U409 ( .B(n526), .A(n527), .S(n1190), .Y(n525) );
  MUX2X1 U410 ( .B(n529), .A(n530), .S(n1190), .Y(n528) );
  MUX2X1 U411 ( .B(n532), .A(n533), .S(n1190), .Y(n531) );
  MUX2X1 U412 ( .B(n535), .A(n536), .S(n1190), .Y(n534) );
  MUX2X1 U413 ( .B(n538), .A(n539), .S(n1175), .Y(n537) );
  MUX2X1 U414 ( .B(n541), .A(n542), .S(n1190), .Y(n540) );
  MUX2X1 U415 ( .B(n544), .A(n545), .S(n1190), .Y(n543) );
  MUX2X1 U416 ( .B(n547), .A(n548), .S(n1190), .Y(n546) );
  MUX2X1 U417 ( .B(n550), .A(n551), .S(n1190), .Y(n549) );
  MUX2X1 U418 ( .B(n553), .A(n554), .S(n1174), .Y(n552) );
  MUX2X1 U419 ( .B(n556), .A(n557), .S(n1191), .Y(n555) );
  MUX2X1 U420 ( .B(n559), .A(n560), .S(n1191), .Y(n558) );
  MUX2X1 U421 ( .B(n562), .A(n563), .S(n1191), .Y(n561) );
  MUX2X1 U422 ( .B(n565), .A(n566), .S(n1191), .Y(n564) );
  MUX2X1 U423 ( .B(n568), .A(n569), .S(n1174), .Y(n567) );
  MUX2X1 U424 ( .B(n571), .A(n572), .S(n1191), .Y(n570) );
  MUX2X1 U425 ( .B(n574), .A(n575), .S(n1191), .Y(n573) );
  MUX2X1 U426 ( .B(n577), .A(n578), .S(n1191), .Y(n576) );
  MUX2X1 U427 ( .B(n580), .A(n581), .S(n1191), .Y(n579) );
  MUX2X1 U428 ( .B(n583), .A(n584), .S(n1174), .Y(n582) );
  MUX2X1 U429 ( .B(n586), .A(n587), .S(n1191), .Y(n585) );
  MUX2X1 U430 ( .B(n589), .A(n590), .S(n1191), .Y(n588) );
  MUX2X1 U431 ( .B(n592), .A(n593), .S(n1191), .Y(n591) );
  MUX2X1 U432 ( .B(n595), .A(n596), .S(n1191), .Y(n594) );
  MUX2X1 U433 ( .B(n598), .A(n599), .S(n1174), .Y(n597) );
  MUX2X1 U434 ( .B(n601), .A(n602), .S(n1192), .Y(n600) );
  MUX2X1 U435 ( .B(n604), .A(n605), .S(n1192), .Y(n603) );
  MUX2X1 U436 ( .B(n607), .A(n608), .S(n1192), .Y(n606) );
  MUX2X1 U437 ( .B(n610), .A(n611), .S(n1192), .Y(n609) );
  MUX2X1 U438 ( .B(n613), .A(n614), .S(n1174), .Y(n612) );
  MUX2X1 U439 ( .B(n616), .A(n617), .S(n1192), .Y(n615) );
  MUX2X1 U440 ( .B(n619), .A(n620), .S(n1192), .Y(n618) );
  MUX2X1 U441 ( .B(n622), .A(n623), .S(n1192), .Y(n621) );
  MUX2X1 U442 ( .B(n625), .A(n626), .S(n1192), .Y(n624) );
  MUX2X1 U443 ( .B(n628), .A(n629), .S(n1175), .Y(n627) );
  MUX2X1 U444 ( .B(n631), .A(n632), .S(n1192), .Y(n630) );
  MUX2X1 U445 ( .B(n634), .A(n635), .S(n1192), .Y(n633) );
  MUX2X1 U446 ( .B(n637), .A(n638), .S(n1192), .Y(n636) );
  MUX2X1 U447 ( .B(n640), .A(n641), .S(n1192), .Y(n639) );
  MUX2X1 U448 ( .B(n643), .A(n644), .S(n1175), .Y(n642) );
  MUX2X1 U449 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n1206), .Y(n166) );
  MUX2X1 U450 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n1205), .Y(n165) );
  MUX2X1 U451 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n1207), .Y(n169) );
  MUX2X1 U452 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n1199), .Y(n168) );
  MUX2X1 U453 ( .B(n167), .A(n164), .S(n1179), .Y(n178) );
  MUX2X1 U454 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n1208), .Y(n172) );
  MUX2X1 U455 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n1202), .Y(n171) );
  MUX2X1 U456 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n1201), .Y(n175) );
  MUX2X1 U457 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n1200), .Y(n174) );
  MUX2X1 U458 ( .B(n173), .A(n170), .S(n1179), .Y(n177) );
  MUX2X1 U459 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n1199), .Y(n181) );
  MUX2X1 U460 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n1206), .Y(n180) );
  MUX2X1 U461 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n1197), .Y(n184) );
  MUX2X1 U462 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n1199), .Y(n183) );
  MUX2X1 U463 ( .B(n182), .A(n179), .S(n1179), .Y(n193) );
  MUX2X1 U464 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n1198), .Y(n187) );
  MUX2X1 U465 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n1209), .Y(n186) );
  MUX2X1 U466 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n1207), .Y(n190) );
  MUX2X1 U467 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n1206), .Y(n189) );
  MUX2X1 U468 ( .B(n188), .A(n185), .S(n1179), .Y(n192) );
  MUX2X1 U469 ( .B(n191), .A(n176), .S(n1173), .Y(n645) );
  MUX2X1 U470 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n1196), .Y(n196) );
  MUX2X1 U471 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n1196), .Y(n195) );
  MUX2X1 U472 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n1196), .Y(n199) );
  MUX2X1 U473 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n1196), .Y(n198) );
  MUX2X1 U474 ( .B(n197), .A(n194), .S(n1179), .Y(n208) );
  MUX2X1 U475 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n1196), .Y(n202) );
  MUX2X1 U476 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n1196), .Y(n201) );
  MUX2X1 U477 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n1196), .Y(n205) );
  MUX2X1 U478 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n1196), .Y(n204) );
  MUX2X1 U479 ( .B(n203), .A(n200), .S(n1179), .Y(n207) );
  MUX2X1 U480 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n1196), .Y(n211) );
  MUX2X1 U481 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n1196), .Y(n210) );
  MUX2X1 U482 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n1196), .Y(n215) );
  MUX2X1 U483 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n1196), .Y(n213) );
  MUX2X1 U484 ( .B(n212), .A(n209), .S(n1179), .Y(n224) );
  MUX2X1 U485 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n1201), .Y(n218) );
  MUX2X1 U486 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n1197), .Y(n217) );
  MUX2X1 U487 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n1209), .Y(n221) );
  MUX2X1 U488 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n1200), .Y(n220) );
  MUX2X1 U489 ( .B(n219), .A(n216), .S(n1179), .Y(n223) );
  MUX2X1 U490 ( .B(n222), .A(n206), .S(n1173), .Y(n646) );
  MUX2X1 U491 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n1199), .Y(n227) );
  MUX2X1 U492 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n1207), .Y(n226) );
  MUX2X1 U493 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n1200), .Y(n230) );
  MUX2X1 U494 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n1209), .Y(n229) );
  MUX2X1 U495 ( .B(n228), .A(n225), .S(n1179), .Y(n239) );
  MUX2X1 U496 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n1211), .Y(n233) );
  MUX2X1 U497 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n1210), .Y(n232) );
  MUX2X1 U498 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n1207), .Y(n236) );
  MUX2X1 U499 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n1197), .Y(n235) );
  MUX2X1 U500 ( .B(n234), .A(n231), .S(n1179), .Y(n238) );
  MUX2X1 U501 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n1209), .Y(n242) );
  MUX2X1 U502 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n1204), .Y(n241) );
  MUX2X1 U503 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n1209), .Y(n245) );
  MUX2X1 U504 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n1198), .Y(n244) );
  MUX2X1 U505 ( .B(n243), .A(n240), .S(n1179), .Y(n254) );
  MUX2X1 U506 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n1208), .Y(n248) );
  MUX2X1 U507 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n1205), .Y(n247) );
  MUX2X1 U508 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n1209), .Y(n251) );
  MUX2X1 U509 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n1202), .Y(n250) );
  MUX2X1 U510 ( .B(n249), .A(n246), .S(n1179), .Y(n253) );
  MUX2X1 U511 ( .B(n252), .A(n237), .S(n1173), .Y(n647) );
  MUX2X1 U512 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n1207), .Y(n257) );
  MUX2X1 U513 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n1203), .Y(n256) );
  MUX2X1 U514 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n1209), .Y(n260) );
  MUX2X1 U515 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n1206), .Y(n259) );
  MUX2X1 U516 ( .B(n258), .A(n255), .S(n1178), .Y(n269) );
  MUX2X1 U517 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n1197), .Y(n263) );
  MUX2X1 U518 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n1197), .Y(n262) );
  MUX2X1 U519 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n1197), .Y(n266) );
  MUX2X1 U520 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n1197), .Y(n265) );
  MUX2X1 U521 ( .B(n264), .A(n261), .S(n1178), .Y(n268) );
  MUX2X1 U522 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n1197), .Y(n272) );
  MUX2X1 U523 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n1197), .Y(n271) );
  MUX2X1 U524 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n1197), .Y(n275) );
  MUX2X1 U525 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n1197), .Y(n274) );
  MUX2X1 U526 ( .B(n273), .A(n270), .S(n1178), .Y(n284) );
  MUX2X1 U527 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n1197), .Y(n278) );
  MUX2X1 U528 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n1197), .Y(n277) );
  MUX2X1 U529 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n1197), .Y(n281) );
  MUX2X1 U530 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n1197), .Y(n280) );
  MUX2X1 U531 ( .B(n279), .A(n276), .S(n1178), .Y(n283) );
  MUX2X1 U532 ( .B(n282), .A(n267), .S(n1173), .Y(n648) );
  MUX2X1 U533 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n1198), .Y(n287) );
  MUX2X1 U534 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n1198), .Y(n286) );
  MUX2X1 U535 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n1198), .Y(n290) );
  MUX2X1 U536 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n1198), .Y(n289) );
  MUX2X1 U537 ( .B(n288), .A(n285), .S(n1178), .Y(n299) );
  MUX2X1 U538 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n1198), .Y(n293) );
  MUX2X1 U539 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n1198), .Y(n292) );
  MUX2X1 U540 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n1198), .Y(n296) );
  MUX2X1 U541 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n1198), .Y(n295) );
  MUX2X1 U542 ( .B(n294), .A(n291), .S(n1178), .Y(n298) );
  MUX2X1 U543 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n1198), .Y(n302) );
  MUX2X1 U544 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n1198), .Y(n301) );
  MUX2X1 U545 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n1198), .Y(n305) );
  MUX2X1 U546 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n1198), .Y(n304) );
  MUX2X1 U547 ( .B(n303), .A(n300), .S(n1178), .Y(n314) );
  MUX2X1 U548 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n1199), .Y(n308) );
  MUX2X1 U549 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n1199), .Y(n307) );
  MUX2X1 U550 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n1199), .Y(n311) );
  MUX2X1 U551 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n1199), .Y(n310) );
  MUX2X1 U552 ( .B(n309), .A(n306), .S(n1178), .Y(n313) );
  MUX2X1 U553 ( .B(n312), .A(n297), .S(n1173), .Y(n649) );
  MUX2X1 U554 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n1199), .Y(n317) );
  MUX2X1 U555 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n1199), .Y(n316) );
  MUX2X1 U556 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n1199), .Y(n320) );
  MUX2X1 U557 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n1199), .Y(n319) );
  MUX2X1 U558 ( .B(n318), .A(n315), .S(n1178), .Y(n329) );
  MUX2X1 U559 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n1199), .Y(n323) );
  MUX2X1 U560 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n1199), .Y(n322) );
  MUX2X1 U561 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n1199), .Y(n326) );
  MUX2X1 U562 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n1199), .Y(n325) );
  MUX2X1 U563 ( .B(n324), .A(n321), .S(n1178), .Y(n328) );
  MUX2X1 U564 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n1206), .Y(n332) );
  MUX2X1 U565 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n1198), .Y(n331) );
  MUX2X1 U566 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n1209), .Y(n335) );
  MUX2X1 U567 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n1209), .Y(n334) );
  MUX2X1 U568 ( .B(n333), .A(n330), .S(n1178), .Y(n344) );
  MUX2X1 U569 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n1209), .Y(n338) );
  MUX2X1 U570 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n1200), .Y(n337) );
  MUX2X1 U571 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n1196), .Y(n341) );
  MUX2X1 U572 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n1201), .Y(n340) );
  MUX2X1 U573 ( .B(n339), .A(n336), .S(n1178), .Y(n343) );
  MUX2X1 U574 ( .B(n342), .A(n327), .S(n1173), .Y(n650) );
  MUX2X1 U575 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n1201), .Y(n347) );
  MUX2X1 U576 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n1206), .Y(n346) );
  MUX2X1 U577 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n1208), .Y(n350) );
  MUX2X1 U578 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n1207), .Y(n349) );
  MUX2X1 U579 ( .B(n348), .A(n345), .S(n1178), .Y(n359) );
  MUX2X1 U580 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n1200), .Y(n353) );
  MUX2X1 U581 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n1200), .Y(n352) );
  MUX2X1 U582 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n1200), .Y(n356) );
  MUX2X1 U583 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n1200), .Y(n355) );
  MUX2X1 U584 ( .B(n354), .A(n351), .S(n1179), .Y(n358) );
  MUX2X1 U585 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n1200), .Y(n362) );
  MUX2X1 U586 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n1200), .Y(n361) );
  MUX2X1 U587 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n1200), .Y(n365) );
  MUX2X1 U588 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n1200), .Y(n364) );
  MUX2X1 U589 ( .B(n363), .A(n360), .S(n1178), .Y(n374) );
  MUX2X1 U590 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n1200), .Y(n368) );
  MUX2X1 U591 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n1200), .Y(n367) );
  MUX2X1 U592 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n1200), .Y(n371) );
  MUX2X1 U593 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n1200), .Y(n370) );
  MUX2X1 U594 ( .B(n369), .A(n366), .S(n1179), .Y(n373) );
  MUX2X1 U595 ( .B(n372), .A(n357), .S(n1173), .Y(n1163) );
  MUX2X1 U596 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n1201), .Y(n377) );
  MUX2X1 U597 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n1201), .Y(n376) );
  MUX2X1 U598 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n1201), .Y(n380) );
  MUX2X1 U599 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n1201), .Y(n379) );
  MUX2X1 U600 ( .B(n378), .A(n375), .S(n1179), .Y(n389) );
  MUX2X1 U601 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n1201), .Y(n383) );
  MUX2X1 U602 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n1201), .Y(n382) );
  MUX2X1 U603 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n1201), .Y(n386) );
  MUX2X1 U604 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n1201), .Y(n385) );
  MUX2X1 U605 ( .B(n384), .A(n381), .S(n1178), .Y(n388) );
  MUX2X1 U606 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n1201), .Y(n392) );
  MUX2X1 U607 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n1201), .Y(n391) );
  MUX2X1 U608 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n1201), .Y(n395) );
  MUX2X1 U609 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n1201), .Y(n394) );
  MUX2X1 U610 ( .B(n393), .A(n390), .S(n1179), .Y(n404) );
  MUX2X1 U611 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n1202), .Y(n398) );
  MUX2X1 U612 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n1202), .Y(n397) );
  MUX2X1 U613 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n1202), .Y(n401) );
  MUX2X1 U614 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n1202), .Y(n400) );
  MUX2X1 U615 ( .B(n399), .A(n396), .S(n1178), .Y(n403) );
  MUX2X1 U616 ( .B(n402), .A(n387), .S(n1173), .Y(n1164) );
  MUX2X1 U617 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n1202), .Y(n407) );
  MUX2X1 U618 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n1202), .Y(n406) );
  MUX2X1 U619 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n1202), .Y(n410) );
  MUX2X1 U620 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n1202), .Y(n409) );
  MUX2X1 U621 ( .B(n408), .A(n405), .S(n1179), .Y(n419) );
  MUX2X1 U622 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n1202), .Y(n413) );
  MUX2X1 U623 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n1202), .Y(n412) );
  MUX2X1 U624 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n1202), .Y(n416) );
  MUX2X1 U625 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n1202), .Y(n415) );
  MUX2X1 U626 ( .B(n414), .A(n411), .S(n1178), .Y(n418) );
  MUX2X1 U627 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n1203), .Y(n422) );
  MUX2X1 U628 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n1203), .Y(n421) );
  MUX2X1 U629 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n1203), .Y(n425) );
  MUX2X1 U630 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n1203), .Y(n424) );
  MUX2X1 U631 ( .B(n423), .A(n420), .S(n1178), .Y(n434) );
  MUX2X1 U632 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n1203), .Y(n428) );
  MUX2X1 U633 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n1203), .Y(n427) );
  MUX2X1 U634 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n1203), .Y(n431) );
  MUX2X1 U635 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n1203), .Y(n430) );
  MUX2X1 U636 ( .B(n429), .A(n426), .S(n1178), .Y(n433) );
  MUX2X1 U637 ( .B(n432), .A(n417), .S(n1173), .Y(n1165) );
  MUX2X1 U638 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n1203), .Y(n437) );
  MUX2X1 U639 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n1203), .Y(n436) );
  MUX2X1 U640 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n1203), .Y(n440) );
  MUX2X1 U641 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n1203), .Y(n439) );
  MUX2X1 U642 ( .B(n438), .A(n435), .S(n1177), .Y(n449) );
  MUX2X1 U643 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n1204), .Y(n443) );
  MUX2X1 U644 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n1204), .Y(n442) );
  MUX2X1 U645 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n1204), .Y(n446) );
  MUX2X1 U646 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n1204), .Y(n445) );
  MUX2X1 U647 ( .B(n444), .A(n441), .S(n1177), .Y(n448) );
  MUX2X1 U648 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n1204), .Y(n452) );
  MUX2X1 U649 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n1204), .Y(n451) );
  MUX2X1 U650 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n1204), .Y(n455) );
  MUX2X1 U651 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n1204), .Y(n454) );
  MUX2X1 U652 ( .B(n453), .A(n450), .S(n1177), .Y(n464) );
  MUX2X1 U653 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n1204), .Y(n458) );
  MUX2X1 U654 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n1204), .Y(n457) );
  MUX2X1 U655 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n1204), .Y(n461) );
  MUX2X1 U656 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n1204), .Y(n460) );
  MUX2X1 U657 ( .B(n459), .A(n456), .S(n1177), .Y(n463) );
  MUX2X1 U658 ( .B(n462), .A(n447), .S(n1173), .Y(n1166) );
  MUX2X1 U659 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n1205), .Y(n467) );
  MUX2X1 U660 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n1205), .Y(n466) );
  MUX2X1 U661 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n1205), .Y(n470) );
  MUX2X1 U662 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n1205), .Y(n469) );
  MUX2X1 U663 ( .B(n468), .A(n465), .S(n1177), .Y(n479) );
  MUX2X1 U664 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n1205), .Y(n473) );
  MUX2X1 U665 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n1205), .Y(n472) );
  MUX2X1 U666 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n1205), .Y(n476) );
  MUX2X1 U667 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n1205), .Y(n475) );
  MUX2X1 U668 ( .B(n474), .A(n471), .S(n1177), .Y(n478) );
  MUX2X1 U669 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n1205), .Y(n482) );
  MUX2X1 U670 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n1205), .Y(n481) );
  MUX2X1 U671 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n1205), .Y(n485) );
  MUX2X1 U672 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n1205), .Y(n484) );
  MUX2X1 U673 ( .B(n483), .A(n480), .S(n1177), .Y(n494) );
  MUX2X1 U674 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n1206), .Y(n488) );
  MUX2X1 U675 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n1206), .Y(n487) );
  MUX2X1 U676 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n1206), .Y(n491) );
  MUX2X1 U677 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n1206), .Y(n490) );
  MUX2X1 U678 ( .B(n489), .A(n486), .S(n1177), .Y(n493) );
  MUX2X1 U679 ( .B(n492), .A(n477), .S(n1173), .Y(n1167) );
  MUX2X1 U680 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n1206), .Y(n497) );
  MUX2X1 U681 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n1206), .Y(n496) );
  MUX2X1 U682 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n1206), .Y(n500) );
  MUX2X1 U683 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n1206), .Y(n499) );
  MUX2X1 U684 ( .B(n498), .A(n495), .S(n1177), .Y(n509) );
  MUX2X1 U685 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n1206), .Y(n503) );
  MUX2X1 U686 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n1206), .Y(n502) );
  MUX2X1 U687 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n1206), .Y(n506) );
  MUX2X1 U688 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n1206), .Y(n505) );
  MUX2X1 U689 ( .B(n504), .A(n501), .S(n1177), .Y(n508) );
  MUX2X1 U690 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n1207), .Y(n512) );
  MUX2X1 U691 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n1207), .Y(n511) );
  MUX2X1 U692 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n1207), .Y(n515) );
  MUX2X1 U693 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n1207), .Y(n514) );
  MUX2X1 U694 ( .B(n513), .A(n510), .S(n1177), .Y(n524) );
  MUX2X1 U695 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n1207), .Y(n518) );
  MUX2X1 U696 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n1207), .Y(n517) );
  MUX2X1 U697 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n1207), .Y(n521) );
  MUX2X1 U698 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n1207), .Y(n520) );
  MUX2X1 U699 ( .B(n519), .A(n516), .S(n1177), .Y(n523) );
  MUX2X1 U700 ( .B(n522), .A(n507), .S(n1173), .Y(n1168) );
  MUX2X1 U701 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n1207), .Y(n527) );
  MUX2X1 U702 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n1207), .Y(n526) );
  MUX2X1 U703 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n1207), .Y(n530) );
  MUX2X1 U704 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n1207), .Y(n529) );
  MUX2X1 U705 ( .B(n528), .A(n525), .S(n1176), .Y(n539) );
  MUX2X1 U706 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n1208), .Y(n533) );
  MUX2X1 U707 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n1208), .Y(n532) );
  MUX2X1 U708 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n1208), .Y(n536) );
  MUX2X1 U709 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n1208), .Y(n535) );
  MUX2X1 U710 ( .B(n534), .A(n531), .S(n1176), .Y(n538) );
  MUX2X1 U711 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n1208), .Y(n542) );
  MUX2X1 U712 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n1208), .Y(n541) );
  MUX2X1 U713 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n1208), .Y(n545) );
  MUX2X1 U714 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n1208), .Y(n544) );
  MUX2X1 U715 ( .B(n543), .A(n540), .S(n1176), .Y(n554) );
  MUX2X1 U716 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n1208), .Y(n548) );
  MUX2X1 U717 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n1208), .Y(n547) );
  MUX2X1 U718 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n1208), .Y(n551) );
  MUX2X1 U719 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n1208), .Y(n550) );
  MUX2X1 U720 ( .B(n549), .A(n546), .S(n1176), .Y(n553) );
  MUX2X1 U721 ( .B(n552), .A(n537), .S(n1173), .Y(n1169) );
  MUX2X1 U722 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n1209), .Y(n557) );
  MUX2X1 U723 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n1209), .Y(n556) );
  MUX2X1 U724 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n1209), .Y(n560) );
  MUX2X1 U725 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n1209), .Y(n559) );
  MUX2X1 U726 ( .B(n558), .A(n555), .S(n1176), .Y(n569) );
  MUX2X1 U727 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n1209), .Y(n563) );
  MUX2X1 U728 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n1209), .Y(n562) );
  MUX2X1 U729 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n1209), .Y(n566) );
  MUX2X1 U730 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n1209), .Y(n565) );
  MUX2X1 U731 ( .B(n564), .A(n561), .S(n1176), .Y(n568) );
  MUX2X1 U732 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n1209), .Y(n572) );
  MUX2X1 U733 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n1209), .Y(n571) );
  MUX2X1 U734 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n1209), .Y(n575) );
  MUX2X1 U735 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n1209), .Y(n574) );
  MUX2X1 U736 ( .B(n573), .A(n570), .S(n1176), .Y(n584) );
  MUX2X1 U737 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n1210), .Y(n578) );
  MUX2X1 U738 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n1210), .Y(n577) );
  MUX2X1 U739 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n1210), .Y(n581) );
  MUX2X1 U740 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n1210), .Y(n580) );
  MUX2X1 U741 ( .B(n579), .A(n576), .S(n1176), .Y(n583) );
  MUX2X1 U742 ( .B(n582), .A(n567), .S(n1173), .Y(n1170) );
  MUX2X1 U743 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n1210), .Y(n587) );
  MUX2X1 U744 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n1210), .Y(n586) );
  MUX2X1 U745 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n1210), .Y(n590) );
  MUX2X1 U746 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n1210), .Y(n589) );
  MUX2X1 U747 ( .B(n588), .A(n585), .S(n1176), .Y(n599) );
  MUX2X1 U748 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n1210), .Y(n593) );
  MUX2X1 U749 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n1210), .Y(n592) );
  MUX2X1 U750 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n1210), .Y(n596) );
  MUX2X1 U751 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n1210), .Y(n595) );
  MUX2X1 U752 ( .B(n594), .A(n591), .S(n1176), .Y(n598) );
  MUX2X1 U753 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n1211), .Y(n602) );
  MUX2X1 U754 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n1211), .Y(n601) );
  MUX2X1 U755 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n1211), .Y(n605) );
  MUX2X1 U756 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n1211), .Y(n604) );
  MUX2X1 U757 ( .B(n603), .A(n600), .S(n1176), .Y(n614) );
  MUX2X1 U758 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n1211), .Y(n608) );
  MUX2X1 U759 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n1211), .Y(n607) );
  MUX2X1 U760 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n1211), .Y(n611) );
  MUX2X1 U761 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n1211), .Y(n610) );
  MUX2X1 U762 ( .B(n609), .A(n606), .S(n1176), .Y(n613) );
  MUX2X1 U763 ( .B(n612), .A(n597), .S(n1173), .Y(n1171) );
  MUX2X1 U764 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n1211), .Y(n617) );
  MUX2X1 U765 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n1211), .Y(n616) );
  MUX2X1 U766 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n1211), .Y(n620) );
  MUX2X1 U767 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n1211), .Y(n619) );
  MUX2X1 U768 ( .B(n618), .A(n615), .S(n1177), .Y(n629) );
  MUX2X1 U769 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n1202), .Y(n623) );
  MUX2X1 U770 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n1202), .Y(n622) );
  MUX2X1 U771 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n1208), .Y(n626) );
  MUX2X1 U772 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n1199), .Y(n625) );
  MUX2X1 U773 ( .B(n624), .A(n621), .S(n1176), .Y(n628) );
  MUX2X1 U774 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n1198), .Y(n632) );
  MUX2X1 U775 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n1202), .Y(n631) );
  MUX2X1 U776 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n1212), .Y(n635) );
  MUX2X1 U777 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n1208), .Y(n634) );
  MUX2X1 U778 ( .B(n633), .A(n630), .S(n1177), .Y(n644) );
  MUX2X1 U779 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n1199), .Y(n638) );
  MUX2X1 U780 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n1196), .Y(n637) );
  MUX2X1 U781 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n1212), .Y(n641) );
  MUX2X1 U782 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n1197), .Y(n640) );
  MUX2X1 U783 ( .B(n639), .A(n636), .S(n1176), .Y(n643) );
  MUX2X1 U784 ( .B(n642), .A(n627), .S(n1173), .Y(n1172) );
  INVX8 U785 ( .A(n1296), .Y(n1212) );
  INVX1 U786 ( .A(N12), .Y(n1299) );
  INVX1 U787 ( .A(N11), .Y(n1298) );
  INVX8 U788 ( .A(n1270), .Y(n1267) );
  INVX8 U789 ( .A(n1270), .Y(n1268) );
  INVX8 U790 ( .A(n1270), .Y(n1269) );
  INVX8 U791 ( .A(n76), .Y(n1271) );
  INVX8 U792 ( .A(n76), .Y(n1272) );
  INVX8 U793 ( .A(n77), .Y(n1273) );
  INVX8 U794 ( .A(n78), .Y(n1274) );
  INVX8 U795 ( .A(n79), .Y(n1275) );
  INVX8 U796 ( .A(n80), .Y(n1276) );
  INVX8 U797 ( .A(n80), .Y(n1277) );
  INVX8 U798 ( .A(n81), .Y(n1278) );
  INVX8 U799 ( .A(n82), .Y(n1279) );
  INVX8 U800 ( .A(n83), .Y(n1280) );
  INVX8 U801 ( .A(n84), .Y(n1281) );
  INVX8 U802 ( .A(n84), .Y(n1282) );
  INVX8 U803 ( .A(n85), .Y(n1283) );
  INVX8 U804 ( .A(n86), .Y(n1284) );
  INVX8 U805 ( .A(n87), .Y(n1285) );
  INVX8 U806 ( .A(n87), .Y(n1286) );
  INVX8 U807 ( .A(n88), .Y(n1287) );
  INVX8 U808 ( .A(n88), .Y(n1288) );
  INVX8 U809 ( .A(n89), .Y(n1289) );
  INVX8 U810 ( .A(n89), .Y(n1290) );
  INVX8 U811 ( .A(n90), .Y(n1291) );
  INVX8 U812 ( .A(n90), .Y(n1292) );
  INVX8 U813 ( .A(n91), .Y(n1293) );
  INVX8 U814 ( .A(n91), .Y(n1294) );
  OR2X2 U815 ( .A(write), .B(rst), .Y(n1303) );
  AND2X2 U816 ( .A(N32), .B(n3), .Y(\data_out<0> ) );
  AND2X2 U817 ( .A(n4), .B(N31), .Y(\data_out<1> ) );
  AND2X2 U818 ( .A(N30), .B(n1304), .Y(\data_out<2> ) );
  AND2X2 U819 ( .A(n4), .B(N29), .Y(\data_out<3> ) );
  AND2X2 U820 ( .A(n4), .B(N28), .Y(\data_out<4> ) );
  AND2X2 U821 ( .A(n4), .B(N27), .Y(\data_out<5> ) );
  AND2X2 U822 ( .A(n4), .B(N26), .Y(\data_out<6> ) );
  AND2X2 U823 ( .A(N25), .B(n3), .Y(\data_out<7> ) );
  AND2X2 U824 ( .A(N24), .B(n4), .Y(\data_out<8> ) );
  AND2X2 U825 ( .A(N23), .B(n1304), .Y(\data_out<9> ) );
  AND2X2 U826 ( .A(N22), .B(n3), .Y(\data_out<10> ) );
  AND2X2 U827 ( .A(N21), .B(n4), .Y(\data_out<11> ) );
  AND2X2 U828 ( .A(N20), .B(n4), .Y(\data_out<12> ) );
  AND2X2 U829 ( .A(N19), .B(n1304), .Y(\data_out<13> ) );
  AND2X2 U830 ( .A(N18), .B(n3), .Y(\data_out<14> ) );
  AND2X2 U831 ( .A(N17), .B(n3), .Y(\data_out<15> ) );
  NAND2X1 U832 ( .A(\mem<31><0> ), .B(n1213), .Y(n1305) );
  OAI21X1 U833 ( .A(n97), .B(n1271), .C(n1305), .Y(n2343) );
  NAND2X1 U834 ( .A(\mem<31><1> ), .B(n1213), .Y(n1306) );
  OAI21X1 U835 ( .A(n1273), .B(n97), .C(n1306), .Y(n2342) );
  NAND2X1 U836 ( .A(\mem<31><2> ), .B(n1213), .Y(n1307) );
  OAI21X1 U837 ( .A(n1274), .B(n97), .C(n1307), .Y(n2341) );
  NAND2X1 U838 ( .A(\mem<31><3> ), .B(n1213), .Y(n1308) );
  OAI21X1 U839 ( .A(n1275), .B(n97), .C(n1308), .Y(n2340) );
  NAND2X1 U840 ( .A(\mem<31><4> ), .B(n1213), .Y(n1309) );
  OAI21X1 U841 ( .A(n1277), .B(n97), .C(n1309), .Y(n2339) );
  NAND2X1 U842 ( .A(\mem<31><5> ), .B(n1213), .Y(n1310) );
  OAI21X1 U843 ( .A(n1278), .B(n97), .C(n1310), .Y(n2338) );
  NAND2X1 U844 ( .A(\mem<31><6> ), .B(n1213), .Y(n1311) );
  OAI21X1 U845 ( .A(n1279), .B(n97), .C(n1311), .Y(n2337) );
  NAND2X1 U846 ( .A(\mem<31><7> ), .B(n1213), .Y(n1312) );
  OAI21X1 U847 ( .A(n1280), .B(n97), .C(n1312), .Y(n2336) );
  NAND2X1 U848 ( .A(\mem<31><8> ), .B(n1214), .Y(n1313) );
  OAI21X1 U849 ( .A(n1282), .B(n97), .C(n1313), .Y(n2335) );
  NAND2X1 U850 ( .A(\mem<31><9> ), .B(n1214), .Y(n1314) );
  OAI21X1 U851 ( .A(n1283), .B(n97), .C(n1314), .Y(n2334) );
  NAND2X1 U852 ( .A(\mem<31><10> ), .B(n1214), .Y(n1315) );
  OAI21X1 U853 ( .A(n1284), .B(n97), .C(n1315), .Y(n2333) );
  NAND2X1 U854 ( .A(\mem<31><11> ), .B(n1214), .Y(n1316) );
  OAI21X1 U855 ( .A(n1286), .B(n97), .C(n1316), .Y(n2332) );
  NAND2X1 U856 ( .A(\mem<31><12> ), .B(n1214), .Y(n1317) );
  OAI21X1 U857 ( .A(n1288), .B(n97), .C(n1317), .Y(n2331) );
  NAND2X1 U858 ( .A(\mem<31><13> ), .B(n1214), .Y(n1318) );
  OAI21X1 U859 ( .A(n1290), .B(n97), .C(n1318), .Y(n2330) );
  NAND2X1 U860 ( .A(\mem<31><14> ), .B(n1214), .Y(n1319) );
  OAI21X1 U861 ( .A(n1292), .B(n97), .C(n1319), .Y(n2329) );
  NAND2X1 U862 ( .A(\mem<31><15> ), .B(n1214), .Y(n1320) );
  OAI21X1 U863 ( .A(n1294), .B(n97), .C(n1320), .Y(n2328) );
  NAND2X1 U864 ( .A(\mem<30><0> ), .B(n1215), .Y(n1321) );
  OAI21X1 U865 ( .A(n99), .B(n1271), .C(n1321), .Y(n2327) );
  NAND2X1 U866 ( .A(\mem<30><1> ), .B(n1215), .Y(n1322) );
  OAI21X1 U867 ( .A(n99), .B(n1273), .C(n1322), .Y(n2326) );
  NAND2X1 U868 ( .A(\mem<30><2> ), .B(n1215), .Y(n1323) );
  OAI21X1 U869 ( .A(n99), .B(n1274), .C(n1323), .Y(n2325) );
  NAND2X1 U870 ( .A(\mem<30><3> ), .B(n1215), .Y(n1324) );
  OAI21X1 U871 ( .A(n99), .B(n1275), .C(n1324), .Y(n2324) );
  NAND2X1 U872 ( .A(\mem<30><4> ), .B(n1215), .Y(n1325) );
  OAI21X1 U873 ( .A(n99), .B(n1277), .C(n1325), .Y(n2323) );
  NAND2X1 U874 ( .A(\mem<30><5> ), .B(n1215), .Y(n1326) );
  OAI21X1 U875 ( .A(n99), .B(n1278), .C(n1326), .Y(n2322) );
  NAND2X1 U876 ( .A(\mem<30><6> ), .B(n1215), .Y(n1327) );
  OAI21X1 U877 ( .A(n99), .B(n1279), .C(n1327), .Y(n2321) );
  NAND2X1 U878 ( .A(\mem<30><7> ), .B(n1215), .Y(n1328) );
  OAI21X1 U879 ( .A(n99), .B(n1280), .C(n1328), .Y(n2320) );
  NAND2X1 U880 ( .A(\mem<30><8> ), .B(n1216), .Y(n1329) );
  OAI21X1 U881 ( .A(n99), .B(n1281), .C(n1329), .Y(n2319) );
  NAND2X1 U882 ( .A(\mem<30><9> ), .B(n1216), .Y(n1330) );
  OAI21X1 U883 ( .A(n99), .B(n1283), .C(n1330), .Y(n2318) );
  NAND2X1 U884 ( .A(\mem<30><10> ), .B(n1216), .Y(n1331) );
  OAI21X1 U885 ( .A(n99), .B(n1284), .C(n1331), .Y(n2317) );
  NAND2X1 U886 ( .A(\mem<30><11> ), .B(n1216), .Y(n1332) );
  OAI21X1 U887 ( .A(n99), .B(n1285), .C(n1332), .Y(n2316) );
  NAND2X1 U888 ( .A(\mem<30><12> ), .B(n1216), .Y(n1333) );
  OAI21X1 U889 ( .A(n99), .B(n1287), .C(n1333), .Y(n2315) );
  NAND2X1 U890 ( .A(\mem<30><13> ), .B(n1216), .Y(n1334) );
  OAI21X1 U891 ( .A(n99), .B(n1289), .C(n1334), .Y(n2314) );
  NAND2X1 U892 ( .A(\mem<30><14> ), .B(n1216), .Y(n1335) );
  OAI21X1 U893 ( .A(n99), .B(n1291), .C(n1335), .Y(n2313) );
  NAND2X1 U894 ( .A(\mem<30><15> ), .B(n1216), .Y(n1336) );
  OAI21X1 U895 ( .A(n99), .B(n1293), .C(n1336), .Y(n2312) );
  NAND3X1 U896 ( .A(n1196), .B(n1176), .C(n1298), .Y(n1337) );
  NAND2X1 U897 ( .A(\mem<29><0> ), .B(n1217), .Y(n1338) );
  OAI21X1 U898 ( .A(n101), .B(n1271), .C(n1338), .Y(n2311) );
  NAND2X1 U899 ( .A(\mem<29><1> ), .B(n1217), .Y(n1339) );
  OAI21X1 U900 ( .A(n101), .B(n1273), .C(n1339), .Y(n2310) );
  NAND2X1 U901 ( .A(\mem<29><2> ), .B(n1217), .Y(n1340) );
  OAI21X1 U902 ( .A(n101), .B(n1274), .C(n1340), .Y(n2309) );
  NAND2X1 U903 ( .A(\mem<29><3> ), .B(n1217), .Y(n1341) );
  OAI21X1 U904 ( .A(n101), .B(n1275), .C(n1341), .Y(n2308) );
  NAND2X1 U905 ( .A(\mem<29><4> ), .B(n1217), .Y(n1342) );
  OAI21X1 U906 ( .A(n101), .B(n1276), .C(n1342), .Y(n2307) );
  NAND2X1 U907 ( .A(\mem<29><5> ), .B(n1217), .Y(n1343) );
  OAI21X1 U908 ( .A(n101), .B(n1278), .C(n1343), .Y(n2306) );
  NAND2X1 U909 ( .A(\mem<29><6> ), .B(n1217), .Y(n1344) );
  OAI21X1 U910 ( .A(n101), .B(n1279), .C(n1344), .Y(n2305) );
  NAND2X1 U911 ( .A(\mem<29><7> ), .B(n1217), .Y(n1345) );
  OAI21X1 U912 ( .A(n101), .B(n1280), .C(n1345), .Y(n2304) );
  NAND2X1 U913 ( .A(\mem<29><8> ), .B(n1218), .Y(n1346) );
  OAI21X1 U914 ( .A(n101), .B(n1282), .C(n1346), .Y(n2303) );
  NAND2X1 U915 ( .A(\mem<29><9> ), .B(n1218), .Y(n1347) );
  OAI21X1 U916 ( .A(n101), .B(n1283), .C(n1347), .Y(n2302) );
  NAND2X1 U917 ( .A(\mem<29><10> ), .B(n1218), .Y(n1348) );
  OAI21X1 U918 ( .A(n101), .B(n1284), .C(n1348), .Y(n2301) );
  NAND2X1 U919 ( .A(\mem<29><11> ), .B(n1218), .Y(n1349) );
  OAI21X1 U920 ( .A(n101), .B(n1286), .C(n1349), .Y(n2300) );
  NAND2X1 U921 ( .A(\mem<29><12> ), .B(n1218), .Y(n1350) );
  OAI21X1 U922 ( .A(n101), .B(n1288), .C(n1350), .Y(n2299) );
  NAND2X1 U923 ( .A(\mem<29><13> ), .B(n1218), .Y(n1351) );
  OAI21X1 U924 ( .A(n101), .B(n1290), .C(n1351), .Y(n2298) );
  NAND2X1 U925 ( .A(\mem<29><14> ), .B(n1218), .Y(n1352) );
  OAI21X1 U926 ( .A(n101), .B(n1292), .C(n1352), .Y(n2297) );
  NAND2X1 U927 ( .A(\mem<29><15> ), .B(n1218), .Y(n1353) );
  OAI21X1 U928 ( .A(n101), .B(n1294), .C(n1353), .Y(n2296) );
  NAND3X1 U929 ( .A(n1177), .B(n1298), .C(n1296), .Y(n1354) );
  NAND2X1 U930 ( .A(\mem<28><0> ), .B(n1219), .Y(n1355) );
  OAI21X1 U931 ( .A(n103), .B(n1271), .C(n1355), .Y(n2295) );
  NAND2X1 U932 ( .A(\mem<28><1> ), .B(n1219), .Y(n1356) );
  OAI21X1 U933 ( .A(n103), .B(n1273), .C(n1356), .Y(n2294) );
  NAND2X1 U934 ( .A(\mem<28><2> ), .B(n1219), .Y(n1357) );
  OAI21X1 U935 ( .A(n103), .B(n1274), .C(n1357), .Y(n2293) );
  NAND2X1 U936 ( .A(\mem<28><3> ), .B(n1219), .Y(n1358) );
  OAI21X1 U937 ( .A(n103), .B(n1275), .C(n1358), .Y(n2292) );
  NAND2X1 U938 ( .A(\mem<28><4> ), .B(n1219), .Y(n1359) );
  OAI21X1 U939 ( .A(n103), .B(n1277), .C(n1359), .Y(n2291) );
  NAND2X1 U940 ( .A(\mem<28><5> ), .B(n1219), .Y(n1360) );
  OAI21X1 U941 ( .A(n103), .B(n1278), .C(n1360), .Y(n2290) );
  NAND2X1 U942 ( .A(\mem<28><6> ), .B(n1219), .Y(n1361) );
  OAI21X1 U943 ( .A(n103), .B(n1279), .C(n1361), .Y(n2289) );
  NAND2X1 U944 ( .A(\mem<28><7> ), .B(n1219), .Y(n1362) );
  OAI21X1 U945 ( .A(n103), .B(n1280), .C(n1362), .Y(n2288) );
  NAND2X1 U946 ( .A(\mem<28><8> ), .B(n1220), .Y(n1363) );
  OAI21X1 U947 ( .A(n103), .B(n1281), .C(n1363), .Y(n2287) );
  NAND2X1 U948 ( .A(\mem<28><9> ), .B(n1220), .Y(n1364) );
  OAI21X1 U949 ( .A(n103), .B(n1283), .C(n1364), .Y(n2286) );
  NAND2X1 U950 ( .A(\mem<28><10> ), .B(n1220), .Y(n1365) );
  OAI21X1 U951 ( .A(n103), .B(n1284), .C(n1365), .Y(n2285) );
  NAND2X1 U952 ( .A(\mem<28><11> ), .B(n1220), .Y(n1366) );
  OAI21X1 U953 ( .A(n103), .B(n1285), .C(n1366), .Y(n2284) );
  NAND2X1 U954 ( .A(\mem<28><12> ), .B(n1220), .Y(n1367) );
  OAI21X1 U955 ( .A(n103), .B(n1287), .C(n1367), .Y(n2283) );
  NAND2X1 U956 ( .A(\mem<28><13> ), .B(n1220), .Y(n1368) );
  OAI21X1 U957 ( .A(n103), .B(n1289), .C(n1368), .Y(n2282) );
  NAND2X1 U958 ( .A(\mem<28><14> ), .B(n1220), .Y(n1369) );
  OAI21X1 U959 ( .A(n103), .B(n1291), .C(n1369), .Y(n2281) );
  NAND2X1 U960 ( .A(\mem<28><15> ), .B(n1220), .Y(n1370) );
  OAI21X1 U961 ( .A(n103), .B(n1293), .C(n1370), .Y(n2280) );
  NAND3X1 U962 ( .A(n1196), .B(n1297), .C(n1299), .Y(n1371) );
  NAND2X1 U963 ( .A(\mem<27><0> ), .B(n1221), .Y(n1372) );
  OAI21X1 U964 ( .A(n105), .B(n1271), .C(n1372), .Y(n2279) );
  NAND2X1 U965 ( .A(\mem<27><1> ), .B(n1221), .Y(n1373) );
  OAI21X1 U966 ( .A(n105), .B(n1273), .C(n1373), .Y(n2278) );
  NAND2X1 U967 ( .A(\mem<27><2> ), .B(n1221), .Y(n1374) );
  OAI21X1 U968 ( .A(n105), .B(n1274), .C(n1374), .Y(n2277) );
  NAND2X1 U969 ( .A(\mem<27><3> ), .B(n1221), .Y(n1375) );
  OAI21X1 U970 ( .A(n105), .B(n1275), .C(n1375), .Y(n2276) );
  NAND2X1 U971 ( .A(\mem<27><4> ), .B(n1221), .Y(n1376) );
  OAI21X1 U972 ( .A(n105), .B(n1276), .C(n1376), .Y(n2275) );
  NAND2X1 U973 ( .A(\mem<27><5> ), .B(n1221), .Y(n1377) );
  OAI21X1 U974 ( .A(n105), .B(n1278), .C(n1377), .Y(n2274) );
  NAND2X1 U975 ( .A(\mem<27><6> ), .B(n1221), .Y(n1378) );
  OAI21X1 U976 ( .A(n105), .B(n1279), .C(n1378), .Y(n2273) );
  NAND2X1 U977 ( .A(\mem<27><7> ), .B(n1221), .Y(n1379) );
  OAI21X1 U978 ( .A(n105), .B(n1280), .C(n1379), .Y(n2272) );
  NAND2X1 U979 ( .A(\mem<27><8> ), .B(n1222), .Y(n1380) );
  OAI21X1 U980 ( .A(n105), .B(n1282), .C(n1380), .Y(n2271) );
  NAND2X1 U981 ( .A(\mem<27><9> ), .B(n1222), .Y(n1381) );
  OAI21X1 U982 ( .A(n105), .B(n1283), .C(n1381), .Y(n2270) );
  NAND2X1 U983 ( .A(\mem<27><10> ), .B(n1222), .Y(n1382) );
  OAI21X1 U984 ( .A(n105), .B(n1284), .C(n1382), .Y(n2269) );
  NAND2X1 U985 ( .A(\mem<27><11> ), .B(n1222), .Y(n1383) );
  OAI21X1 U986 ( .A(n105), .B(n1286), .C(n1383), .Y(n2268) );
  NAND2X1 U987 ( .A(\mem<27><12> ), .B(n1222), .Y(n1384) );
  OAI21X1 U988 ( .A(n105), .B(n1288), .C(n1384), .Y(n2267) );
  NAND2X1 U989 ( .A(\mem<27><13> ), .B(n1222), .Y(n1385) );
  OAI21X1 U990 ( .A(n105), .B(n1290), .C(n1385), .Y(n2266) );
  NAND2X1 U991 ( .A(\mem<27><14> ), .B(n1222), .Y(n1386) );
  OAI21X1 U992 ( .A(n105), .B(n1292), .C(n1386), .Y(n2265) );
  NAND2X1 U993 ( .A(\mem<27><15> ), .B(n1222), .Y(n1387) );
  OAI21X1 U994 ( .A(n105), .B(n1294), .C(n1387), .Y(n2264) );
  NAND3X1 U995 ( .A(n1299), .B(n1297), .C(n1296), .Y(n1388) );
  NAND2X1 U996 ( .A(\mem<26><0> ), .B(n1223), .Y(n1389) );
  OAI21X1 U997 ( .A(n107), .B(n1271), .C(n1389), .Y(n2263) );
  NAND2X1 U998 ( .A(\mem<26><1> ), .B(n1223), .Y(n1390) );
  OAI21X1 U999 ( .A(n107), .B(n1273), .C(n1390), .Y(n2262) );
  NAND2X1 U1000 ( .A(\mem<26><2> ), .B(n1223), .Y(n1391) );
  OAI21X1 U1001 ( .A(n107), .B(n1274), .C(n1391), .Y(n2261) );
  NAND2X1 U1002 ( .A(\mem<26><3> ), .B(n1223), .Y(n1392) );
  OAI21X1 U1003 ( .A(n107), .B(n1275), .C(n1392), .Y(n2260) );
  NAND2X1 U1004 ( .A(\mem<26><4> ), .B(n1223), .Y(n1393) );
  OAI21X1 U1005 ( .A(n107), .B(n1277), .C(n1393), .Y(n2259) );
  NAND2X1 U1006 ( .A(\mem<26><5> ), .B(n1223), .Y(n1394) );
  OAI21X1 U1007 ( .A(n107), .B(n1278), .C(n1394), .Y(n2258) );
  NAND2X1 U1008 ( .A(\mem<26><6> ), .B(n1223), .Y(n1395) );
  OAI21X1 U1009 ( .A(n107), .B(n1279), .C(n1395), .Y(n2257) );
  NAND2X1 U1010 ( .A(\mem<26><7> ), .B(n1223), .Y(n1396) );
  OAI21X1 U1011 ( .A(n107), .B(n1280), .C(n1396), .Y(n2256) );
  NAND2X1 U1012 ( .A(\mem<26><8> ), .B(n1224), .Y(n1397) );
  OAI21X1 U1013 ( .A(n107), .B(n1281), .C(n1397), .Y(n2255) );
  NAND2X1 U1014 ( .A(\mem<26><9> ), .B(n1224), .Y(n1398) );
  OAI21X1 U1015 ( .A(n107), .B(n1283), .C(n1398), .Y(n2254) );
  NAND2X1 U1016 ( .A(\mem<26><10> ), .B(n1224), .Y(n1399) );
  OAI21X1 U1017 ( .A(n107), .B(n1284), .C(n1399), .Y(n2253) );
  NAND2X1 U1018 ( .A(\mem<26><11> ), .B(n1224), .Y(n1400) );
  OAI21X1 U1019 ( .A(n107), .B(n1285), .C(n1400), .Y(n2252) );
  NAND2X1 U1020 ( .A(\mem<26><12> ), .B(n1224), .Y(n1401) );
  OAI21X1 U1021 ( .A(n107), .B(n1287), .C(n1401), .Y(n2251) );
  NAND2X1 U1022 ( .A(\mem<26><13> ), .B(n1224), .Y(n1402) );
  OAI21X1 U1023 ( .A(n107), .B(n1289), .C(n1402), .Y(n2250) );
  NAND2X1 U1024 ( .A(\mem<26><14> ), .B(n1224), .Y(n1403) );
  OAI21X1 U1025 ( .A(n107), .B(n1291), .C(n1403), .Y(n2249) );
  NAND2X1 U1026 ( .A(\mem<26><15> ), .B(n1224), .Y(n1404) );
  OAI21X1 U1027 ( .A(n107), .B(n1293), .C(n1404), .Y(n2248) );
  NAND3X1 U1028 ( .A(n1196), .B(n1299), .C(n1298), .Y(n1405) );
  NAND2X1 U1029 ( .A(\mem<25><0> ), .B(n1225), .Y(n1406) );
  OAI21X1 U1030 ( .A(n109), .B(n1271), .C(n1406), .Y(n2247) );
  NAND2X1 U1031 ( .A(\mem<25><1> ), .B(n1225), .Y(n1407) );
  OAI21X1 U1032 ( .A(n109), .B(n1273), .C(n1407), .Y(n2246) );
  NAND2X1 U1033 ( .A(\mem<25><2> ), .B(n1225), .Y(n1408) );
  OAI21X1 U1034 ( .A(n109), .B(n1274), .C(n1408), .Y(n2245) );
  NAND2X1 U1035 ( .A(\mem<25><3> ), .B(n1225), .Y(n1409) );
  OAI21X1 U1036 ( .A(n109), .B(n1275), .C(n1409), .Y(n2244) );
  NAND2X1 U1037 ( .A(\mem<25><4> ), .B(n1225), .Y(n1410) );
  OAI21X1 U1038 ( .A(n109), .B(n1276), .C(n1410), .Y(n2243) );
  NAND2X1 U1039 ( .A(\mem<25><5> ), .B(n1225), .Y(n1411) );
  OAI21X1 U1040 ( .A(n109), .B(n1278), .C(n1411), .Y(n2242) );
  NAND2X1 U1041 ( .A(\mem<25><6> ), .B(n1225), .Y(n1412) );
  OAI21X1 U1042 ( .A(n109), .B(n1279), .C(n1412), .Y(n2241) );
  NAND2X1 U1043 ( .A(\mem<25><7> ), .B(n1225), .Y(n1413) );
  OAI21X1 U1044 ( .A(n109), .B(n1280), .C(n1413), .Y(n2240) );
  NAND2X1 U1045 ( .A(\mem<25><8> ), .B(n1226), .Y(n1414) );
  OAI21X1 U1046 ( .A(n109), .B(n1282), .C(n1414), .Y(n2239) );
  NAND2X1 U1047 ( .A(\mem<25><9> ), .B(n1226), .Y(n1415) );
  OAI21X1 U1048 ( .A(n109), .B(n1283), .C(n1415), .Y(n2238) );
  NAND2X1 U1049 ( .A(\mem<25><10> ), .B(n1226), .Y(n1416) );
  OAI21X1 U1050 ( .A(n109), .B(n1284), .C(n1416), .Y(n2237) );
  NAND2X1 U1051 ( .A(\mem<25><11> ), .B(n1226), .Y(n1417) );
  OAI21X1 U1052 ( .A(n109), .B(n1286), .C(n1417), .Y(n2236) );
  NAND2X1 U1053 ( .A(\mem<25><12> ), .B(n1226), .Y(n1418) );
  OAI21X1 U1054 ( .A(n109), .B(n1288), .C(n1418), .Y(n2235) );
  NAND2X1 U1055 ( .A(\mem<25><13> ), .B(n1226), .Y(n1419) );
  OAI21X1 U1056 ( .A(n109), .B(n1290), .C(n1419), .Y(n2234) );
  NAND2X1 U1057 ( .A(\mem<25><14> ), .B(n1226), .Y(n1420) );
  OAI21X1 U1058 ( .A(n109), .B(n1292), .C(n1420), .Y(n2233) );
  NAND2X1 U1059 ( .A(\mem<25><15> ), .B(n1226), .Y(n1421) );
  OAI21X1 U1060 ( .A(n109), .B(n1294), .C(n1421), .Y(n2232) );
  NOR3X1 U1061 ( .A(n1196), .B(n1297), .C(n1176), .Y(n1815) );
  NAND2X1 U1062 ( .A(\mem<24><0> ), .B(n1228), .Y(n1422) );
  OAI21X1 U1063 ( .A(n1227), .B(n1271), .C(n1422), .Y(n2231) );
  NAND2X1 U1064 ( .A(\mem<24><1> ), .B(n1228), .Y(n1423) );
  OAI21X1 U1065 ( .A(n1227), .B(n1273), .C(n1423), .Y(n2230) );
  NAND2X1 U1066 ( .A(\mem<24><2> ), .B(n1228), .Y(n1424) );
  OAI21X1 U1067 ( .A(n1227), .B(n1274), .C(n1424), .Y(n2229) );
  NAND2X1 U1068 ( .A(\mem<24><3> ), .B(n1228), .Y(n1425) );
  OAI21X1 U1069 ( .A(n1227), .B(n1275), .C(n1425), .Y(n2228) );
  NAND2X1 U1070 ( .A(\mem<24><4> ), .B(n1228), .Y(n1426) );
  OAI21X1 U1071 ( .A(n1227), .B(n1276), .C(n1426), .Y(n2227) );
  NAND2X1 U1072 ( .A(\mem<24><5> ), .B(n1228), .Y(n1427) );
  OAI21X1 U1073 ( .A(n1227), .B(n1278), .C(n1427), .Y(n2226) );
  NAND2X1 U1074 ( .A(\mem<24><6> ), .B(n1228), .Y(n1428) );
  OAI21X1 U1075 ( .A(n1227), .B(n1279), .C(n1428), .Y(n2225) );
  NAND2X1 U1076 ( .A(\mem<24><7> ), .B(n1228), .Y(n1429) );
  OAI21X1 U1077 ( .A(n1227), .B(n1280), .C(n1429), .Y(n2224) );
  NAND2X1 U1078 ( .A(\mem<24><8> ), .B(n1229), .Y(n1430) );
  OAI21X1 U1079 ( .A(n1227), .B(n1281), .C(n1430), .Y(n2223) );
  NAND2X1 U1080 ( .A(\mem<24><9> ), .B(n1229), .Y(n1431) );
  OAI21X1 U1081 ( .A(n1227), .B(n1283), .C(n1431), .Y(n2222) );
  NAND2X1 U1082 ( .A(\mem<24><10> ), .B(n1229), .Y(n1432) );
  OAI21X1 U1083 ( .A(n1227), .B(n1284), .C(n1432), .Y(n2221) );
  NAND2X1 U1084 ( .A(\mem<24><11> ), .B(n1229), .Y(n1433) );
  OAI21X1 U1085 ( .A(n1227), .B(n1285), .C(n1433), .Y(n2220) );
  NAND2X1 U1086 ( .A(\mem<24><12> ), .B(n1229), .Y(n1434) );
  OAI21X1 U1087 ( .A(n1227), .B(n1287), .C(n1434), .Y(n2219) );
  NAND2X1 U1088 ( .A(\mem<24><13> ), .B(n1229), .Y(n1435) );
  OAI21X1 U1089 ( .A(n1227), .B(n1289), .C(n1435), .Y(n2218) );
  NAND2X1 U1090 ( .A(\mem<24><14> ), .B(n1229), .Y(n1436) );
  OAI21X1 U1091 ( .A(n1227), .B(n1291), .C(n1436), .Y(n2217) );
  NAND2X1 U1092 ( .A(\mem<24><15> ), .B(n1229), .Y(n1437) );
  OAI21X1 U1093 ( .A(n1227), .B(n1293), .C(n1437), .Y(n2216) );
  NAND2X1 U1094 ( .A(\mem<23><0> ), .B(n1230), .Y(n1438) );
  OAI21X1 U1095 ( .A(n111), .B(n1271), .C(n1438), .Y(n2215) );
  NAND2X1 U1096 ( .A(\mem<23><1> ), .B(n1230), .Y(n1439) );
  OAI21X1 U1097 ( .A(n111), .B(n1273), .C(n1439), .Y(n2214) );
  NAND2X1 U1098 ( .A(\mem<23><2> ), .B(n1230), .Y(n1440) );
  OAI21X1 U1099 ( .A(n111), .B(n1274), .C(n1440), .Y(n2213) );
  NAND2X1 U1100 ( .A(\mem<23><3> ), .B(n1230), .Y(n1441) );
  OAI21X1 U1101 ( .A(n111), .B(n1275), .C(n1441), .Y(n2212) );
  NAND2X1 U1102 ( .A(\mem<23><4> ), .B(n1230), .Y(n1442) );
  OAI21X1 U1103 ( .A(n111), .B(n1277), .C(n1442), .Y(n2211) );
  NAND2X1 U1104 ( .A(\mem<23><5> ), .B(n1230), .Y(n1443) );
  OAI21X1 U1105 ( .A(n111), .B(n1278), .C(n1443), .Y(n2210) );
  NAND2X1 U1106 ( .A(\mem<23><6> ), .B(n1230), .Y(n1444) );
  OAI21X1 U1107 ( .A(n111), .B(n1279), .C(n1444), .Y(n2209) );
  NAND2X1 U1108 ( .A(\mem<23><7> ), .B(n1230), .Y(n1445) );
  OAI21X1 U1109 ( .A(n111), .B(n1280), .C(n1445), .Y(n2208) );
  NAND2X1 U1110 ( .A(\mem<23><8> ), .B(n1231), .Y(n1446) );
  OAI21X1 U1111 ( .A(n111), .B(n1282), .C(n1446), .Y(n2207) );
  NAND2X1 U1112 ( .A(\mem<23><9> ), .B(n1231), .Y(n1447) );
  OAI21X1 U1113 ( .A(n111), .B(n1283), .C(n1447), .Y(n2206) );
  NAND2X1 U1114 ( .A(\mem<23><10> ), .B(n1231), .Y(n1448) );
  OAI21X1 U1115 ( .A(n111), .B(n1284), .C(n1448), .Y(n2205) );
  NAND2X1 U1116 ( .A(\mem<23><11> ), .B(n1231), .Y(n1449) );
  OAI21X1 U1117 ( .A(n111), .B(n1286), .C(n1449), .Y(n2204) );
  NAND2X1 U1118 ( .A(\mem<23><12> ), .B(n1231), .Y(n1450) );
  OAI21X1 U1119 ( .A(n111), .B(n1288), .C(n1450), .Y(n2203) );
  NAND2X1 U1120 ( .A(\mem<23><13> ), .B(n1231), .Y(n1451) );
  OAI21X1 U1121 ( .A(n111), .B(n1290), .C(n1451), .Y(n2202) );
  NAND2X1 U1122 ( .A(\mem<23><14> ), .B(n1231), .Y(n1452) );
  OAI21X1 U1123 ( .A(n111), .B(n1292), .C(n1452), .Y(n2201) );
  NAND2X1 U1124 ( .A(\mem<23><15> ), .B(n1231), .Y(n1453) );
  OAI21X1 U1125 ( .A(n111), .B(n1294), .C(n1453), .Y(n2200) );
  NAND2X1 U1126 ( .A(\mem<22><0> ), .B(n1232), .Y(n1454) );
  OAI21X1 U1127 ( .A(n113), .B(n1271), .C(n1454), .Y(n2199) );
  NAND2X1 U1128 ( .A(\mem<22><1> ), .B(n1232), .Y(n1455) );
  OAI21X1 U1129 ( .A(n113), .B(n1273), .C(n1455), .Y(n2198) );
  NAND2X1 U1130 ( .A(\mem<22><2> ), .B(n1232), .Y(n1456) );
  OAI21X1 U1131 ( .A(n113), .B(n1274), .C(n1456), .Y(n2197) );
  NAND2X1 U1132 ( .A(\mem<22><3> ), .B(n1232), .Y(n1457) );
  OAI21X1 U1133 ( .A(n113), .B(n1275), .C(n1457), .Y(n2196) );
  NAND2X1 U1134 ( .A(\mem<22><4> ), .B(n1232), .Y(n1458) );
  OAI21X1 U1135 ( .A(n113), .B(n1277), .C(n1458), .Y(n2195) );
  NAND2X1 U1136 ( .A(\mem<22><5> ), .B(n1232), .Y(n1459) );
  OAI21X1 U1137 ( .A(n113), .B(n1278), .C(n1459), .Y(n2194) );
  NAND2X1 U1138 ( .A(\mem<22><6> ), .B(n1232), .Y(n1460) );
  OAI21X1 U1139 ( .A(n113), .B(n1279), .C(n1460), .Y(n2193) );
  NAND2X1 U1140 ( .A(\mem<22><7> ), .B(n1232), .Y(n1461) );
  OAI21X1 U1141 ( .A(n113), .B(n1280), .C(n1461), .Y(n2192) );
  NAND2X1 U1142 ( .A(\mem<22><8> ), .B(n1233), .Y(n1462) );
  OAI21X1 U1143 ( .A(n113), .B(n1282), .C(n1462), .Y(n2191) );
  NAND2X1 U1144 ( .A(\mem<22><9> ), .B(n1233), .Y(n1463) );
  OAI21X1 U1145 ( .A(n113), .B(n1283), .C(n1463), .Y(n2190) );
  NAND2X1 U1146 ( .A(\mem<22><10> ), .B(n1233), .Y(n1464) );
  OAI21X1 U1147 ( .A(n113), .B(n1284), .C(n1464), .Y(n2189) );
  NAND2X1 U1148 ( .A(\mem<22><11> ), .B(n1233), .Y(n1465) );
  OAI21X1 U1149 ( .A(n113), .B(n1286), .C(n1465), .Y(n2188) );
  NAND2X1 U1150 ( .A(\mem<22><12> ), .B(n1233), .Y(n1466) );
  OAI21X1 U1151 ( .A(n113), .B(n1288), .C(n1466), .Y(n2187) );
  NAND2X1 U1152 ( .A(\mem<22><13> ), .B(n1233), .Y(n1467) );
  OAI21X1 U1153 ( .A(n113), .B(n1290), .C(n1467), .Y(n2186) );
  NAND2X1 U1154 ( .A(\mem<22><14> ), .B(n1233), .Y(n1468) );
  OAI21X1 U1155 ( .A(n113), .B(n1292), .C(n1468), .Y(n2185) );
  NAND2X1 U1156 ( .A(\mem<22><15> ), .B(n1233), .Y(n1469) );
  OAI21X1 U1157 ( .A(n113), .B(n1294), .C(n1469), .Y(n2184) );
  NAND2X1 U1158 ( .A(\mem<21><0> ), .B(n1234), .Y(n1470) );
  OAI21X1 U1159 ( .A(n115), .B(n1271), .C(n1470), .Y(n2183) );
  NAND2X1 U1160 ( .A(\mem<21><1> ), .B(n1234), .Y(n1471) );
  OAI21X1 U1161 ( .A(n115), .B(n1273), .C(n1471), .Y(n2182) );
  NAND2X1 U1162 ( .A(\mem<21><2> ), .B(n1234), .Y(n1472) );
  OAI21X1 U1163 ( .A(n115), .B(n1274), .C(n1472), .Y(n2181) );
  NAND2X1 U1164 ( .A(\mem<21><3> ), .B(n1234), .Y(n1473) );
  OAI21X1 U1165 ( .A(n115), .B(n1275), .C(n1473), .Y(n2180) );
  NAND2X1 U1166 ( .A(\mem<21><4> ), .B(n1234), .Y(n1474) );
  OAI21X1 U1167 ( .A(n115), .B(n1277), .C(n1474), .Y(n2179) );
  NAND2X1 U1168 ( .A(\mem<21><5> ), .B(n1234), .Y(n1475) );
  OAI21X1 U1169 ( .A(n115), .B(n1278), .C(n1475), .Y(n2178) );
  NAND2X1 U1170 ( .A(\mem<21><6> ), .B(n1234), .Y(n1476) );
  OAI21X1 U1171 ( .A(n115), .B(n1279), .C(n1476), .Y(n2177) );
  NAND2X1 U1172 ( .A(\mem<21><7> ), .B(n1234), .Y(n1477) );
  OAI21X1 U1173 ( .A(n115), .B(n1280), .C(n1477), .Y(n2176) );
  NAND2X1 U1174 ( .A(\mem<21><8> ), .B(n1235), .Y(n1478) );
  OAI21X1 U1175 ( .A(n115), .B(n1282), .C(n1478), .Y(n2175) );
  NAND2X1 U1177 ( .A(\mem<21><9> ), .B(n1235), .Y(n1479) );
  OAI21X1 U1178 ( .A(n115), .B(n1283), .C(n1479), .Y(n2174) );
  NAND2X1 U1179 ( .A(\mem<21><10> ), .B(n1235), .Y(n1480) );
  OAI21X1 U1180 ( .A(n115), .B(n1284), .C(n1480), .Y(n2173) );
  NAND2X1 U1181 ( .A(\mem<21><11> ), .B(n1235), .Y(n1481) );
  OAI21X1 U1182 ( .A(n115), .B(n1286), .C(n1481), .Y(n2172) );
  NAND2X1 U1183 ( .A(\mem<21><12> ), .B(n1235), .Y(n1482) );
  OAI21X1 U1184 ( .A(n115), .B(n1288), .C(n1482), .Y(n2171) );
  NAND2X1 U1185 ( .A(\mem<21><13> ), .B(n1235), .Y(n1483) );
  OAI21X1 U1186 ( .A(n115), .B(n1290), .C(n1483), .Y(n2170) );
  NAND2X1 U1187 ( .A(\mem<21><14> ), .B(n1235), .Y(n1484) );
  OAI21X1 U1188 ( .A(n115), .B(n1292), .C(n1484), .Y(n2169) );
  NAND2X1 U1189 ( .A(\mem<21><15> ), .B(n1235), .Y(n1485) );
  OAI21X1 U1190 ( .A(n115), .B(n1294), .C(n1485), .Y(n2168) );
  NAND2X1 U1191 ( .A(\mem<20><0> ), .B(n1236), .Y(n1486) );
  OAI21X1 U1192 ( .A(n117), .B(n1271), .C(n1486), .Y(n2167) );
  NAND2X1 U1193 ( .A(\mem<20><1> ), .B(n1236), .Y(n1487) );
  OAI21X1 U1194 ( .A(n117), .B(n1273), .C(n1487), .Y(n2166) );
  NAND2X1 U1195 ( .A(\mem<20><2> ), .B(n1236), .Y(n1488) );
  OAI21X1 U1196 ( .A(n117), .B(n1274), .C(n1488), .Y(n2165) );
  NAND2X1 U1197 ( .A(\mem<20><3> ), .B(n1236), .Y(n1489) );
  OAI21X1 U1198 ( .A(n117), .B(n1275), .C(n1489), .Y(n2164) );
  NAND2X1 U1199 ( .A(\mem<20><4> ), .B(n1236), .Y(n1490) );
  OAI21X1 U1200 ( .A(n117), .B(n1277), .C(n1490), .Y(n2163) );
  NAND2X1 U1201 ( .A(\mem<20><5> ), .B(n1236), .Y(n1491) );
  OAI21X1 U1202 ( .A(n117), .B(n1278), .C(n1491), .Y(n2162) );
  NAND2X1 U1203 ( .A(\mem<20><6> ), .B(n1236), .Y(n1492) );
  OAI21X1 U1204 ( .A(n117), .B(n1279), .C(n1492), .Y(n2161) );
  NAND2X1 U1205 ( .A(\mem<20><7> ), .B(n1236), .Y(n1493) );
  OAI21X1 U1206 ( .A(n117), .B(n1280), .C(n1493), .Y(n2160) );
  NAND2X1 U1207 ( .A(\mem<20><8> ), .B(n1237), .Y(n1494) );
  OAI21X1 U1208 ( .A(n117), .B(n1282), .C(n1494), .Y(n2159) );
  NAND2X1 U1209 ( .A(\mem<20><9> ), .B(n1237), .Y(n1495) );
  OAI21X1 U1210 ( .A(n117), .B(n1283), .C(n1495), .Y(n2158) );
  NAND2X1 U1211 ( .A(\mem<20><10> ), .B(n1237), .Y(n1496) );
  OAI21X1 U1212 ( .A(n117), .B(n1284), .C(n1496), .Y(n2157) );
  NAND2X1 U1213 ( .A(\mem<20><11> ), .B(n1237), .Y(n1497) );
  OAI21X1 U1214 ( .A(n117), .B(n1286), .C(n1497), .Y(n2156) );
  NAND2X1 U1215 ( .A(\mem<20><12> ), .B(n1237), .Y(n1498) );
  OAI21X1 U1216 ( .A(n117), .B(n1288), .C(n1498), .Y(n2155) );
  NAND2X1 U1217 ( .A(\mem<20><13> ), .B(n1237), .Y(n1499) );
  OAI21X1 U1218 ( .A(n117), .B(n1290), .C(n1499), .Y(n2154) );
  NAND2X1 U1219 ( .A(\mem<20><14> ), .B(n1237), .Y(n1500) );
  OAI21X1 U1220 ( .A(n117), .B(n1292), .C(n1500), .Y(n2153) );
  NAND2X1 U1221 ( .A(\mem<20><15> ), .B(n1237), .Y(n1501) );
  OAI21X1 U1222 ( .A(n117), .B(n1294), .C(n1501), .Y(n2152) );
  NAND2X1 U1223 ( .A(\mem<19><0> ), .B(n1238), .Y(n1502) );
  OAI21X1 U1224 ( .A(n119), .B(n1272), .C(n1502), .Y(n2151) );
  NAND2X1 U1225 ( .A(\mem<19><1> ), .B(n1238), .Y(n1503) );
  OAI21X1 U1226 ( .A(n119), .B(n1273), .C(n1503), .Y(n2150) );
  NAND2X1 U1227 ( .A(\mem<19><2> ), .B(n1238), .Y(n1504) );
  OAI21X1 U1228 ( .A(n119), .B(n1274), .C(n1504), .Y(n2149) );
  NAND2X1 U1229 ( .A(\mem<19><3> ), .B(n1238), .Y(n1505) );
  OAI21X1 U1230 ( .A(n119), .B(n1275), .C(n1505), .Y(n2148) );
  NAND2X1 U1231 ( .A(\mem<19><4> ), .B(n1238), .Y(n1506) );
  OAI21X1 U1232 ( .A(n119), .B(n1277), .C(n1506), .Y(n2147) );
  NAND2X1 U1233 ( .A(\mem<19><5> ), .B(n1238), .Y(n1507) );
  OAI21X1 U1234 ( .A(n119), .B(n1278), .C(n1507), .Y(n2146) );
  NAND2X1 U1235 ( .A(\mem<19><6> ), .B(n1238), .Y(n1508) );
  OAI21X1 U1236 ( .A(n119), .B(n1279), .C(n1508), .Y(n2145) );
  NAND2X1 U1237 ( .A(\mem<19><7> ), .B(n1238), .Y(n1509) );
  OAI21X1 U1238 ( .A(n119), .B(n1280), .C(n1509), .Y(n2144) );
  NAND2X1 U1239 ( .A(\mem<19><8> ), .B(n1239), .Y(n1510) );
  OAI21X1 U1240 ( .A(n119), .B(n1282), .C(n1510), .Y(n2143) );
  NAND2X1 U1241 ( .A(\mem<19><9> ), .B(n1239), .Y(n1511) );
  OAI21X1 U1242 ( .A(n119), .B(n1283), .C(n1511), .Y(n2142) );
  NAND2X1 U1243 ( .A(\mem<19><10> ), .B(n1239), .Y(n1512) );
  OAI21X1 U1244 ( .A(n119), .B(n1284), .C(n1512), .Y(n2141) );
  NAND2X1 U1245 ( .A(\mem<19><11> ), .B(n1239), .Y(n1513) );
  OAI21X1 U1246 ( .A(n119), .B(n1286), .C(n1513), .Y(n2140) );
  NAND2X1 U1247 ( .A(\mem<19><12> ), .B(n1239), .Y(n1514) );
  OAI21X1 U1248 ( .A(n119), .B(n1288), .C(n1514), .Y(n2139) );
  NAND2X1 U1249 ( .A(\mem<19><13> ), .B(n1239), .Y(n1515) );
  OAI21X1 U1250 ( .A(n119), .B(n1290), .C(n1515), .Y(n2138) );
  NAND2X1 U1251 ( .A(\mem<19><14> ), .B(n1239), .Y(n1516) );
  OAI21X1 U1252 ( .A(n119), .B(n1292), .C(n1516), .Y(n2137) );
  NAND2X1 U1253 ( .A(\mem<19><15> ), .B(n1239), .Y(n1517) );
  OAI21X1 U1254 ( .A(n119), .B(n1294), .C(n1517), .Y(n2136) );
  NAND2X1 U1255 ( .A(\mem<18><0> ), .B(n1240), .Y(n1518) );
  OAI21X1 U1256 ( .A(n121), .B(n1272), .C(n1518), .Y(n2135) );
  NAND2X1 U1257 ( .A(\mem<18><1> ), .B(n1240), .Y(n1519) );
  OAI21X1 U1258 ( .A(n121), .B(n1273), .C(n1519), .Y(n2134) );
  NAND2X1 U1259 ( .A(\mem<18><2> ), .B(n1240), .Y(n1520) );
  OAI21X1 U1260 ( .A(n121), .B(n1274), .C(n1520), .Y(n2133) );
  NAND2X1 U1261 ( .A(\mem<18><3> ), .B(n1240), .Y(n1521) );
  OAI21X1 U1262 ( .A(n121), .B(n1275), .C(n1521), .Y(n2132) );
  NAND2X1 U1263 ( .A(\mem<18><4> ), .B(n1240), .Y(n1522) );
  OAI21X1 U1264 ( .A(n121), .B(n1277), .C(n1522), .Y(n2131) );
  NAND2X1 U1265 ( .A(\mem<18><5> ), .B(n1240), .Y(n1523) );
  OAI21X1 U1266 ( .A(n121), .B(n1278), .C(n1523), .Y(n2130) );
  NAND2X1 U1267 ( .A(\mem<18><6> ), .B(n1240), .Y(n1524) );
  OAI21X1 U1268 ( .A(n121), .B(n1279), .C(n1524), .Y(n2129) );
  NAND2X1 U1269 ( .A(\mem<18><7> ), .B(n1240), .Y(n1525) );
  OAI21X1 U1270 ( .A(n121), .B(n1280), .C(n1525), .Y(n2128) );
  NAND2X1 U1271 ( .A(\mem<18><8> ), .B(n1241), .Y(n1526) );
  OAI21X1 U1272 ( .A(n121), .B(n1282), .C(n1526), .Y(n2127) );
  NAND2X1 U1273 ( .A(\mem<18><9> ), .B(n1241), .Y(n1527) );
  OAI21X1 U1274 ( .A(n121), .B(n1283), .C(n1527), .Y(n2126) );
  NAND2X1 U1275 ( .A(\mem<18><10> ), .B(n1241), .Y(n1528) );
  OAI21X1 U1276 ( .A(n121), .B(n1284), .C(n1528), .Y(n2125) );
  NAND2X1 U1277 ( .A(\mem<18><11> ), .B(n1241), .Y(n1529) );
  OAI21X1 U1278 ( .A(n121), .B(n1286), .C(n1529), .Y(n2124) );
  NAND2X1 U1279 ( .A(\mem<18><12> ), .B(n1241), .Y(n1530) );
  OAI21X1 U1280 ( .A(n121), .B(n1288), .C(n1530), .Y(n2123) );
  NAND2X1 U1281 ( .A(\mem<18><13> ), .B(n1241), .Y(n1531) );
  OAI21X1 U1282 ( .A(n121), .B(n1290), .C(n1531), .Y(n2122) );
  NAND2X1 U1283 ( .A(\mem<18><14> ), .B(n1241), .Y(n1532) );
  OAI21X1 U1284 ( .A(n121), .B(n1292), .C(n1532), .Y(n2121) );
  NAND2X1 U1285 ( .A(\mem<18><15> ), .B(n1241), .Y(n1533) );
  OAI21X1 U1286 ( .A(n121), .B(n1294), .C(n1533), .Y(n2120) );
  NAND2X1 U1287 ( .A(\mem<17><0> ), .B(n1242), .Y(n1534) );
  OAI21X1 U1288 ( .A(n123), .B(n1272), .C(n1534), .Y(n2119) );
  NAND2X1 U1289 ( .A(\mem<17><1> ), .B(n1242), .Y(n1535) );
  OAI21X1 U1290 ( .A(n123), .B(n1273), .C(n1535), .Y(n2118) );
  NAND2X1 U1291 ( .A(\mem<17><2> ), .B(n1242), .Y(n1536) );
  OAI21X1 U1292 ( .A(n123), .B(n1274), .C(n1536), .Y(n2117) );
  NAND2X1 U1293 ( .A(\mem<17><3> ), .B(n1242), .Y(n1537) );
  OAI21X1 U1294 ( .A(n123), .B(n1275), .C(n1537), .Y(n2116) );
  NAND2X1 U1295 ( .A(\mem<17><4> ), .B(n1242), .Y(n1538) );
  OAI21X1 U1296 ( .A(n123), .B(n1277), .C(n1538), .Y(n2115) );
  NAND2X1 U1297 ( .A(\mem<17><5> ), .B(n1242), .Y(n1539) );
  OAI21X1 U1298 ( .A(n123), .B(n1278), .C(n1539), .Y(n2114) );
  NAND2X1 U1299 ( .A(\mem<17><6> ), .B(n1242), .Y(n1540) );
  OAI21X1 U1300 ( .A(n123), .B(n1279), .C(n1540), .Y(n2113) );
  NAND2X1 U1301 ( .A(\mem<17><7> ), .B(n1242), .Y(n1541) );
  OAI21X1 U1302 ( .A(n123), .B(n1280), .C(n1541), .Y(n2112) );
  NAND2X1 U1303 ( .A(\mem<17><8> ), .B(n1243), .Y(n1542) );
  OAI21X1 U1304 ( .A(n123), .B(n1282), .C(n1542), .Y(n2111) );
  NAND2X1 U1305 ( .A(\mem<17><9> ), .B(n1243), .Y(n1543) );
  OAI21X1 U1306 ( .A(n123), .B(n1283), .C(n1543), .Y(n2110) );
  NAND2X1 U1307 ( .A(\mem<17><10> ), .B(n1243), .Y(n1544) );
  OAI21X1 U1308 ( .A(n123), .B(n1284), .C(n1544), .Y(n2109) );
  NAND2X1 U1309 ( .A(\mem<17><11> ), .B(n1243), .Y(n1545) );
  OAI21X1 U1310 ( .A(n123), .B(n1286), .C(n1545), .Y(n2108) );
  NAND2X1 U1311 ( .A(\mem<17><12> ), .B(n1243), .Y(n1546) );
  OAI21X1 U1312 ( .A(n123), .B(n1288), .C(n1546), .Y(n2107) );
  NAND2X1 U1313 ( .A(\mem<17><13> ), .B(n1243), .Y(n1547) );
  OAI21X1 U1314 ( .A(n123), .B(n1290), .C(n1547), .Y(n2106) );
  NAND2X1 U1315 ( .A(\mem<17><14> ), .B(n1243), .Y(n1548) );
  OAI21X1 U1316 ( .A(n123), .B(n1292), .C(n1548), .Y(n2105) );
  NAND2X1 U1317 ( .A(\mem<17><15> ), .B(n1243), .Y(n1549) );
  OAI21X1 U1318 ( .A(n123), .B(n1294), .C(n1549), .Y(n2104) );
  NAND2X1 U1319 ( .A(\mem<16><0> ), .B(n1245), .Y(n1550) );
  OAI21X1 U1320 ( .A(n1244), .B(n1272), .C(n1550), .Y(n2103) );
  NAND2X1 U1321 ( .A(\mem<16><1> ), .B(n1245), .Y(n1551) );
  OAI21X1 U1322 ( .A(n1244), .B(n1273), .C(n1551), .Y(n2102) );
  NAND2X1 U1323 ( .A(\mem<16><2> ), .B(n1245), .Y(n1552) );
  OAI21X1 U1324 ( .A(n1244), .B(n1274), .C(n1552), .Y(n2101) );
  NAND2X1 U1325 ( .A(\mem<16><3> ), .B(n1245), .Y(n1553) );
  OAI21X1 U1326 ( .A(n1244), .B(n1275), .C(n1553), .Y(n2100) );
  NAND2X1 U1327 ( .A(\mem<16><4> ), .B(n1245), .Y(n1554) );
  OAI21X1 U1328 ( .A(n1244), .B(n1277), .C(n1554), .Y(n2099) );
  NAND2X1 U1329 ( .A(\mem<16><5> ), .B(n1245), .Y(n1555) );
  OAI21X1 U1330 ( .A(n1244), .B(n1278), .C(n1555), .Y(n2098) );
  NAND2X1 U1331 ( .A(\mem<16><6> ), .B(n1245), .Y(n1556) );
  OAI21X1 U1332 ( .A(n1244), .B(n1279), .C(n1556), .Y(n2097) );
  NAND2X1 U1333 ( .A(\mem<16><7> ), .B(n1245), .Y(n1557) );
  OAI21X1 U1334 ( .A(n1244), .B(n1280), .C(n1557), .Y(n2096) );
  NAND2X1 U1335 ( .A(\mem<16><8> ), .B(n1246), .Y(n1558) );
  OAI21X1 U1336 ( .A(n1244), .B(n1282), .C(n1558), .Y(n2095) );
  NAND2X1 U1337 ( .A(\mem<16><9> ), .B(n1246), .Y(n1559) );
  OAI21X1 U1338 ( .A(n1244), .B(n1283), .C(n1559), .Y(n2094) );
  NAND2X1 U1339 ( .A(\mem<16><10> ), .B(n1246), .Y(n1560) );
  OAI21X1 U1340 ( .A(n1244), .B(n1284), .C(n1560), .Y(n2093) );
  NAND2X1 U1341 ( .A(\mem<16><11> ), .B(n1246), .Y(n1561) );
  OAI21X1 U1342 ( .A(n1244), .B(n1286), .C(n1561), .Y(n2092) );
  NAND2X1 U1343 ( .A(\mem<16><12> ), .B(n1246), .Y(n1562) );
  OAI21X1 U1344 ( .A(n1244), .B(n1288), .C(n1562), .Y(n2091) );
  NAND2X1 U1345 ( .A(\mem<16><13> ), .B(n1246), .Y(n1563) );
  OAI21X1 U1346 ( .A(n1244), .B(n1290), .C(n1563), .Y(n2090) );
  NAND2X1 U1347 ( .A(\mem<16><14> ), .B(n1246), .Y(n1564) );
  OAI21X1 U1348 ( .A(n1244), .B(n1292), .C(n1564), .Y(n2089) );
  NAND2X1 U1349 ( .A(\mem<16><15> ), .B(n1246), .Y(n1565) );
  OAI21X1 U1350 ( .A(n1244), .B(n1294), .C(n1565), .Y(n2088) );
  NAND3X1 U1351 ( .A(n1175), .B(n2344), .C(n1302), .Y(n1566) );
  NAND2X1 U1352 ( .A(\mem<15><0> ), .B(n1247), .Y(n1567) );
  OAI21X1 U1353 ( .A(n125), .B(n1272), .C(n1567), .Y(n2087) );
  NAND2X1 U1354 ( .A(\mem<15><1> ), .B(n1247), .Y(n1568) );
  OAI21X1 U1355 ( .A(n125), .B(n1273), .C(n1568), .Y(n2086) );
  NAND2X1 U1356 ( .A(\mem<15><2> ), .B(n1247), .Y(n1569) );
  OAI21X1 U1357 ( .A(n125), .B(n1274), .C(n1569), .Y(n2085) );
  NAND2X1 U1358 ( .A(\mem<15><3> ), .B(n1247), .Y(n1570) );
  OAI21X1 U1359 ( .A(n125), .B(n1275), .C(n1570), .Y(n2084) );
  NAND2X1 U1360 ( .A(\mem<15><4> ), .B(n1247), .Y(n1571) );
  OAI21X1 U1361 ( .A(n125), .B(n1277), .C(n1571), .Y(n2083) );
  NAND2X1 U1362 ( .A(\mem<15><5> ), .B(n1247), .Y(n1572) );
  OAI21X1 U1363 ( .A(n125), .B(n1278), .C(n1572), .Y(n2082) );
  NAND2X1 U1364 ( .A(\mem<15><6> ), .B(n1247), .Y(n1573) );
  OAI21X1 U1365 ( .A(n125), .B(n1279), .C(n1573), .Y(n2081) );
  NAND2X1 U1366 ( .A(\mem<15><7> ), .B(n1247), .Y(n1574) );
  OAI21X1 U1367 ( .A(n125), .B(n1280), .C(n1574), .Y(n2080) );
  NAND2X1 U1368 ( .A(\mem<15><8> ), .B(n1248), .Y(n1575) );
  OAI21X1 U1369 ( .A(n125), .B(n1282), .C(n1575), .Y(n2079) );
  NAND2X1 U1370 ( .A(\mem<15><9> ), .B(n1248), .Y(n1576) );
  OAI21X1 U1371 ( .A(n125), .B(n1283), .C(n1576), .Y(n2078) );
  NAND2X1 U1372 ( .A(\mem<15><10> ), .B(n1248), .Y(n1577) );
  OAI21X1 U1373 ( .A(n125), .B(n1284), .C(n1577), .Y(n2077) );
  NAND2X1 U1374 ( .A(\mem<15><11> ), .B(n1248), .Y(n1578) );
  OAI21X1 U1375 ( .A(n125), .B(n1286), .C(n1578), .Y(n2076) );
  NAND2X1 U1376 ( .A(\mem<15><12> ), .B(n1248), .Y(n1579) );
  OAI21X1 U1377 ( .A(n125), .B(n1288), .C(n1579), .Y(n2075) );
  NAND2X1 U1378 ( .A(\mem<15><13> ), .B(n1248), .Y(n1580) );
  OAI21X1 U1379 ( .A(n125), .B(n1290), .C(n1580), .Y(n2074) );
  NAND2X1 U1380 ( .A(\mem<15><14> ), .B(n1248), .Y(n1581) );
  OAI21X1 U1381 ( .A(n125), .B(n1292), .C(n1581), .Y(n2073) );
  NAND2X1 U1382 ( .A(\mem<15><15> ), .B(n1248), .Y(n1582) );
  OAI21X1 U1383 ( .A(n125), .B(n1294), .C(n1582), .Y(n2072) );
  NAND2X1 U1384 ( .A(\mem<14><0> ), .B(n1249), .Y(n1583) );
  OAI21X1 U1385 ( .A(n127), .B(n1272), .C(n1583), .Y(n2071) );
  NAND2X1 U1386 ( .A(\mem<14><1> ), .B(n1249), .Y(n1584) );
  OAI21X1 U1387 ( .A(n127), .B(n1273), .C(n1584), .Y(n2070) );
  NAND2X1 U1388 ( .A(\mem<14><2> ), .B(n1249), .Y(n1585) );
  OAI21X1 U1389 ( .A(n127), .B(n1274), .C(n1585), .Y(n2069) );
  NAND2X1 U1390 ( .A(\mem<14><3> ), .B(n1249), .Y(n1586) );
  OAI21X1 U1391 ( .A(n127), .B(n1275), .C(n1586), .Y(n2068) );
  NAND2X1 U1392 ( .A(\mem<14><4> ), .B(n1249), .Y(n1587) );
  OAI21X1 U1393 ( .A(n127), .B(n1277), .C(n1587), .Y(n2067) );
  NAND2X1 U1394 ( .A(\mem<14><5> ), .B(n1249), .Y(n1588) );
  OAI21X1 U1395 ( .A(n127), .B(n1278), .C(n1588), .Y(n2066) );
  NAND2X1 U1396 ( .A(\mem<14><6> ), .B(n1249), .Y(n1589) );
  OAI21X1 U1397 ( .A(n127), .B(n1279), .C(n1589), .Y(n2065) );
  NAND2X1 U1398 ( .A(\mem<14><7> ), .B(n1249), .Y(n1590) );
  OAI21X1 U1399 ( .A(n127), .B(n1280), .C(n1590), .Y(n2064) );
  NAND2X1 U1400 ( .A(\mem<14><8> ), .B(n1250), .Y(n1591) );
  OAI21X1 U1401 ( .A(n127), .B(n1282), .C(n1591), .Y(n2063) );
  NAND2X1 U1402 ( .A(\mem<14><9> ), .B(n1250), .Y(n1592) );
  OAI21X1 U1403 ( .A(n127), .B(n1283), .C(n1592), .Y(n2062) );
  NAND2X1 U1404 ( .A(\mem<14><10> ), .B(n1250), .Y(n1593) );
  OAI21X1 U1405 ( .A(n127), .B(n1284), .C(n1593), .Y(n2061) );
  NAND2X1 U1406 ( .A(\mem<14><11> ), .B(n1250), .Y(n1594) );
  OAI21X1 U1407 ( .A(n127), .B(n1286), .C(n1594), .Y(n2060) );
  NAND2X1 U1408 ( .A(\mem<14><12> ), .B(n1250), .Y(n1595) );
  OAI21X1 U1409 ( .A(n127), .B(n1288), .C(n1595), .Y(n2059) );
  NAND2X1 U1410 ( .A(\mem<14><13> ), .B(n1250), .Y(n1596) );
  OAI21X1 U1411 ( .A(n127), .B(n1290), .C(n1596), .Y(n2058) );
  NAND2X1 U1412 ( .A(\mem<14><14> ), .B(n1250), .Y(n1597) );
  OAI21X1 U1413 ( .A(n127), .B(n1292), .C(n1597), .Y(n2057) );
  NAND2X1 U1414 ( .A(\mem<14><15> ), .B(n1250), .Y(n1598) );
  OAI21X1 U1415 ( .A(n127), .B(n1294), .C(n1598), .Y(n2056) );
  NAND2X1 U1416 ( .A(\mem<13><0> ), .B(n1251), .Y(n1599) );
  OAI21X1 U1417 ( .A(n129), .B(n1272), .C(n1599), .Y(n2055) );
  NAND2X1 U1418 ( .A(\mem<13><1> ), .B(n1251), .Y(n1600) );
  OAI21X1 U1419 ( .A(n129), .B(n1273), .C(n1600), .Y(n2054) );
  NAND2X1 U1420 ( .A(\mem<13><2> ), .B(n1251), .Y(n1601) );
  OAI21X1 U1421 ( .A(n129), .B(n1274), .C(n1601), .Y(n2053) );
  NAND2X1 U1422 ( .A(\mem<13><3> ), .B(n1251), .Y(n1602) );
  OAI21X1 U1423 ( .A(n129), .B(n1275), .C(n1602), .Y(n2052) );
  NAND2X1 U1424 ( .A(\mem<13><4> ), .B(n1251), .Y(n1603) );
  OAI21X1 U1425 ( .A(n129), .B(n1277), .C(n1603), .Y(n2051) );
  NAND2X1 U1426 ( .A(\mem<13><5> ), .B(n1251), .Y(n1604) );
  OAI21X1 U1427 ( .A(n129), .B(n1278), .C(n1604), .Y(n2050) );
  NAND2X1 U1428 ( .A(\mem<13><6> ), .B(n1251), .Y(n1605) );
  OAI21X1 U1429 ( .A(n129), .B(n1279), .C(n1605), .Y(n2049) );
  NAND2X1 U1430 ( .A(\mem<13><7> ), .B(n1251), .Y(n1606) );
  OAI21X1 U1431 ( .A(n129), .B(n1280), .C(n1606), .Y(n2048) );
  NAND2X1 U1432 ( .A(\mem<13><8> ), .B(n1252), .Y(n1607) );
  OAI21X1 U1433 ( .A(n129), .B(n1282), .C(n1607), .Y(n2047) );
  NAND2X1 U1434 ( .A(\mem<13><9> ), .B(n1252), .Y(n1608) );
  OAI21X1 U1435 ( .A(n129), .B(n1283), .C(n1608), .Y(n2046) );
  NAND2X1 U1436 ( .A(\mem<13><10> ), .B(n1252), .Y(n1609) );
  OAI21X1 U1437 ( .A(n129), .B(n1284), .C(n1609), .Y(n2045) );
  NAND2X1 U1438 ( .A(\mem<13><11> ), .B(n1252), .Y(n1610) );
  OAI21X1 U1439 ( .A(n129), .B(n1286), .C(n1610), .Y(n2044) );
  NAND2X1 U1440 ( .A(\mem<13><12> ), .B(n1252), .Y(n1611) );
  OAI21X1 U1441 ( .A(n129), .B(n1288), .C(n1611), .Y(n2043) );
  NAND2X1 U1442 ( .A(\mem<13><13> ), .B(n1252), .Y(n1612) );
  OAI21X1 U1443 ( .A(n129), .B(n1290), .C(n1612), .Y(n2042) );
  NAND2X1 U1444 ( .A(\mem<13><14> ), .B(n1252), .Y(n1613) );
  OAI21X1 U1445 ( .A(n129), .B(n1292), .C(n1613), .Y(n2041) );
  NAND2X1 U1446 ( .A(\mem<13><15> ), .B(n1252), .Y(n1614) );
  OAI21X1 U1447 ( .A(n129), .B(n1294), .C(n1614), .Y(n2040) );
  NAND2X1 U1448 ( .A(\mem<12><0> ), .B(n1253), .Y(n1615) );
  OAI21X1 U1449 ( .A(n131), .B(n1272), .C(n1615), .Y(n2039) );
  NAND2X1 U1450 ( .A(\mem<12><1> ), .B(n1253), .Y(n1616) );
  OAI21X1 U1451 ( .A(n131), .B(n1273), .C(n1616), .Y(n2038) );
  NAND2X1 U1452 ( .A(\mem<12><2> ), .B(n1253), .Y(n1617) );
  OAI21X1 U1453 ( .A(n131), .B(n1274), .C(n1617), .Y(n2037) );
  NAND2X1 U1454 ( .A(\mem<12><3> ), .B(n1253), .Y(n1618) );
  OAI21X1 U1455 ( .A(n131), .B(n1275), .C(n1618), .Y(n2036) );
  NAND2X1 U1456 ( .A(\mem<12><4> ), .B(n1253), .Y(n1619) );
  OAI21X1 U1457 ( .A(n131), .B(n1277), .C(n1619), .Y(n2035) );
  NAND2X1 U1458 ( .A(\mem<12><5> ), .B(n1253), .Y(n1620) );
  OAI21X1 U1459 ( .A(n131), .B(n1278), .C(n1620), .Y(n2034) );
  NAND2X1 U1460 ( .A(\mem<12><6> ), .B(n1253), .Y(n1621) );
  OAI21X1 U1461 ( .A(n131), .B(n1279), .C(n1621), .Y(n2033) );
  NAND2X1 U1462 ( .A(\mem<12><7> ), .B(n1253), .Y(n1622) );
  OAI21X1 U1463 ( .A(n131), .B(n1280), .C(n1622), .Y(n2032) );
  NAND2X1 U1464 ( .A(\mem<12><8> ), .B(n1254), .Y(n1623) );
  OAI21X1 U1465 ( .A(n131), .B(n1282), .C(n1623), .Y(n2031) );
  NAND2X1 U1466 ( .A(\mem<12><9> ), .B(n1254), .Y(n1624) );
  OAI21X1 U1467 ( .A(n131), .B(n1283), .C(n1624), .Y(n2030) );
  NAND2X1 U1468 ( .A(\mem<12><10> ), .B(n1254), .Y(n1625) );
  OAI21X1 U1469 ( .A(n131), .B(n1284), .C(n1625), .Y(n2029) );
  NAND2X1 U1470 ( .A(\mem<12><11> ), .B(n1254), .Y(n1626) );
  OAI21X1 U1471 ( .A(n131), .B(n1286), .C(n1626), .Y(n2028) );
  NAND2X1 U1472 ( .A(\mem<12><12> ), .B(n1254), .Y(n1627) );
  OAI21X1 U1473 ( .A(n131), .B(n1288), .C(n1627), .Y(n2027) );
  NAND2X1 U1474 ( .A(\mem<12><13> ), .B(n1254), .Y(n1628) );
  OAI21X1 U1475 ( .A(n131), .B(n1290), .C(n1628), .Y(n2026) );
  NAND2X1 U1476 ( .A(\mem<12><14> ), .B(n1254), .Y(n1629) );
  OAI21X1 U1477 ( .A(n131), .B(n1292), .C(n1629), .Y(n2025) );
  NAND2X1 U1478 ( .A(\mem<12><15> ), .B(n1254), .Y(n1630) );
  OAI21X1 U1479 ( .A(n131), .B(n1294), .C(n1630), .Y(n2024) );
  NAND2X1 U1480 ( .A(\mem<11><0> ), .B(n1255), .Y(n1631) );
  OAI21X1 U1481 ( .A(n133), .B(n1272), .C(n1631), .Y(n2023) );
  NAND2X1 U1482 ( .A(\mem<11><1> ), .B(n1255), .Y(n1632) );
  OAI21X1 U1483 ( .A(n133), .B(n1273), .C(n1632), .Y(n2022) );
  NAND2X1 U1484 ( .A(\mem<11><2> ), .B(n1255), .Y(n1633) );
  OAI21X1 U1485 ( .A(n133), .B(n1274), .C(n1633), .Y(n2021) );
  NAND2X1 U1486 ( .A(\mem<11><3> ), .B(n1255), .Y(n1634) );
  OAI21X1 U1487 ( .A(n133), .B(n1275), .C(n1634), .Y(n2020) );
  NAND2X1 U1488 ( .A(\mem<11><4> ), .B(n1255), .Y(n1635) );
  OAI21X1 U1489 ( .A(n133), .B(n1276), .C(n1635), .Y(n2019) );
  NAND2X1 U1490 ( .A(\mem<11><5> ), .B(n1255), .Y(n1636) );
  OAI21X1 U1491 ( .A(n133), .B(n1278), .C(n1636), .Y(n2018) );
  NAND2X1 U1492 ( .A(\mem<11><6> ), .B(n1255), .Y(n1637) );
  OAI21X1 U1493 ( .A(n133), .B(n1279), .C(n1637), .Y(n2017) );
  NAND2X1 U1494 ( .A(\mem<11><7> ), .B(n1255), .Y(n1638) );
  OAI21X1 U1495 ( .A(n133), .B(n1280), .C(n1638), .Y(n2016) );
  NAND2X1 U1496 ( .A(\mem<11><8> ), .B(n1256), .Y(n1639) );
  OAI21X1 U1497 ( .A(n133), .B(n1281), .C(n1639), .Y(n2015) );
  NAND2X1 U1498 ( .A(\mem<11><9> ), .B(n1256), .Y(n1640) );
  OAI21X1 U1499 ( .A(n133), .B(n1283), .C(n1640), .Y(n2014) );
  NAND2X1 U1500 ( .A(\mem<11><10> ), .B(n1256), .Y(n1641) );
  OAI21X1 U1501 ( .A(n133), .B(n1284), .C(n1641), .Y(n2013) );
  NAND2X1 U1502 ( .A(\mem<11><11> ), .B(n1256), .Y(n1642) );
  OAI21X1 U1503 ( .A(n133), .B(n1285), .C(n1642), .Y(n2012) );
  NAND2X1 U1504 ( .A(\mem<11><12> ), .B(n1256), .Y(n1643) );
  OAI21X1 U1505 ( .A(n133), .B(n1287), .C(n1643), .Y(n2011) );
  NAND2X1 U1506 ( .A(\mem<11><13> ), .B(n1256), .Y(n1644) );
  OAI21X1 U1507 ( .A(n133), .B(n1289), .C(n1644), .Y(n2010) );
  NAND2X1 U1508 ( .A(\mem<11><14> ), .B(n1256), .Y(n1645) );
  OAI21X1 U1509 ( .A(n133), .B(n1291), .C(n1645), .Y(n2009) );
  NAND2X1 U1510 ( .A(\mem<11><15> ), .B(n1256), .Y(n1646) );
  OAI21X1 U1511 ( .A(n133), .B(n1293), .C(n1646), .Y(n2008) );
  NAND2X1 U1512 ( .A(\mem<10><0> ), .B(n1257), .Y(n1647) );
  OAI21X1 U1513 ( .A(n135), .B(n1272), .C(n1647), .Y(n2007) );
  NAND2X1 U1514 ( .A(\mem<10><1> ), .B(n1257), .Y(n1648) );
  OAI21X1 U1515 ( .A(n135), .B(n1273), .C(n1648), .Y(n2006) );
  NAND2X1 U1516 ( .A(\mem<10><2> ), .B(n1257), .Y(n1649) );
  OAI21X1 U1517 ( .A(n135), .B(n1274), .C(n1649), .Y(n2005) );
  NAND2X1 U1518 ( .A(\mem<10><3> ), .B(n1257), .Y(n1650) );
  OAI21X1 U1519 ( .A(n135), .B(n1275), .C(n1650), .Y(n2004) );
  NAND2X1 U1520 ( .A(\mem<10><4> ), .B(n1257), .Y(n1651) );
  OAI21X1 U1521 ( .A(n135), .B(n1276), .C(n1651), .Y(n2003) );
  NAND2X1 U1522 ( .A(\mem<10><5> ), .B(n1257), .Y(n1652) );
  OAI21X1 U1523 ( .A(n135), .B(n1278), .C(n1652), .Y(n2002) );
  NAND2X1 U1524 ( .A(\mem<10><6> ), .B(n1257), .Y(n1653) );
  OAI21X1 U1525 ( .A(n135), .B(n1279), .C(n1653), .Y(n2001) );
  NAND2X1 U1526 ( .A(\mem<10><7> ), .B(n1257), .Y(n1654) );
  OAI21X1 U1527 ( .A(n135), .B(n1280), .C(n1654), .Y(n2000) );
  NAND2X1 U1528 ( .A(\mem<10><8> ), .B(n1258), .Y(n1655) );
  OAI21X1 U1529 ( .A(n135), .B(n1281), .C(n1655), .Y(n1999) );
  NAND2X1 U1530 ( .A(\mem<10><9> ), .B(n1258), .Y(n1656) );
  OAI21X1 U1531 ( .A(n135), .B(n1283), .C(n1656), .Y(n1998) );
  NAND2X1 U1532 ( .A(\mem<10><10> ), .B(n1258), .Y(n1657) );
  OAI21X1 U1533 ( .A(n135), .B(n1284), .C(n1657), .Y(n1997) );
  NAND2X1 U1534 ( .A(\mem<10><11> ), .B(n1258), .Y(n1658) );
  OAI21X1 U1535 ( .A(n135), .B(n1285), .C(n1658), .Y(n1996) );
  NAND2X1 U1536 ( .A(\mem<10><12> ), .B(n1258), .Y(n1659) );
  OAI21X1 U1537 ( .A(n135), .B(n1287), .C(n1659), .Y(n1995) );
  NAND2X1 U1538 ( .A(\mem<10><13> ), .B(n1258), .Y(n1660) );
  OAI21X1 U1539 ( .A(n135), .B(n1289), .C(n1660), .Y(n1994) );
  NAND2X1 U1540 ( .A(\mem<10><14> ), .B(n1258), .Y(n1661) );
  OAI21X1 U1541 ( .A(n135), .B(n1291), .C(n1661), .Y(n1993) );
  NAND2X1 U1542 ( .A(\mem<10><15> ), .B(n1258), .Y(n1662) );
  OAI21X1 U1543 ( .A(n135), .B(n1293), .C(n1662), .Y(n1992) );
  NAND2X1 U1544 ( .A(\mem<9><0> ), .B(n1259), .Y(n1663) );
  OAI21X1 U1545 ( .A(n137), .B(n1272), .C(n1663), .Y(n1991) );
  NAND2X1 U1546 ( .A(\mem<9><1> ), .B(n1259), .Y(n1664) );
  OAI21X1 U1547 ( .A(n137), .B(n1273), .C(n1664), .Y(n1990) );
  NAND2X1 U1548 ( .A(\mem<9><2> ), .B(n1259), .Y(n1665) );
  OAI21X1 U1549 ( .A(n137), .B(n1274), .C(n1665), .Y(n1989) );
  NAND2X1 U1550 ( .A(\mem<9><3> ), .B(n1259), .Y(n1666) );
  OAI21X1 U1551 ( .A(n137), .B(n1275), .C(n1666), .Y(n1988) );
  NAND2X1 U1552 ( .A(\mem<9><4> ), .B(n1259), .Y(n1667) );
  OAI21X1 U1553 ( .A(n137), .B(n1276), .C(n1667), .Y(n1987) );
  NAND2X1 U1554 ( .A(\mem<9><5> ), .B(n1259), .Y(n1668) );
  OAI21X1 U1555 ( .A(n137), .B(n1278), .C(n1668), .Y(n1986) );
  NAND2X1 U1556 ( .A(\mem<9><6> ), .B(n1259), .Y(n1669) );
  OAI21X1 U1557 ( .A(n137), .B(n1279), .C(n1669), .Y(n1985) );
  NAND2X1 U1558 ( .A(\mem<9><7> ), .B(n1259), .Y(n1670) );
  OAI21X1 U1559 ( .A(n137), .B(n1280), .C(n1670), .Y(n1984) );
  NAND2X1 U1560 ( .A(\mem<9><8> ), .B(n1260), .Y(n1671) );
  OAI21X1 U1561 ( .A(n137), .B(n1281), .C(n1671), .Y(n1983) );
  NAND2X1 U1562 ( .A(\mem<9><9> ), .B(n1260), .Y(n1672) );
  OAI21X1 U1563 ( .A(n137), .B(n1283), .C(n1672), .Y(n1982) );
  NAND2X1 U1564 ( .A(\mem<9><10> ), .B(n1260), .Y(n1673) );
  OAI21X1 U1565 ( .A(n137), .B(n1284), .C(n1673), .Y(n1981) );
  NAND2X1 U1566 ( .A(\mem<9><11> ), .B(n1260), .Y(n1674) );
  OAI21X1 U1567 ( .A(n137), .B(n1285), .C(n1674), .Y(n1980) );
  NAND2X1 U1568 ( .A(\mem<9><12> ), .B(n1260), .Y(n1675) );
  OAI21X1 U1569 ( .A(n137), .B(n1287), .C(n1675), .Y(n1979) );
  NAND2X1 U1570 ( .A(\mem<9><13> ), .B(n1260), .Y(n1676) );
  OAI21X1 U1571 ( .A(n137), .B(n1289), .C(n1676), .Y(n1978) );
  NAND2X1 U1572 ( .A(\mem<9><14> ), .B(n1260), .Y(n1677) );
  OAI21X1 U1573 ( .A(n137), .B(n1291), .C(n1677), .Y(n1977) );
  NAND2X1 U1574 ( .A(\mem<9><15> ), .B(n1260), .Y(n1678) );
  OAI21X1 U1575 ( .A(n137), .B(n1293), .C(n1678), .Y(n1976) );
  NAND2X1 U1576 ( .A(\mem<8><0> ), .B(n1262), .Y(n1680) );
  OAI21X1 U1577 ( .A(n1261), .B(n1272), .C(n1680), .Y(n1975) );
  NAND2X1 U1578 ( .A(\mem<8><1> ), .B(n1262), .Y(n1681) );
  OAI21X1 U1579 ( .A(n1261), .B(n1273), .C(n1681), .Y(n1974) );
  NAND2X1 U1580 ( .A(\mem<8><2> ), .B(n1262), .Y(n1682) );
  OAI21X1 U1581 ( .A(n1261), .B(n1274), .C(n1682), .Y(n1973) );
  NAND2X1 U1582 ( .A(\mem<8><3> ), .B(n1262), .Y(n1683) );
  OAI21X1 U1583 ( .A(n1261), .B(n1275), .C(n1683), .Y(n1972) );
  NAND2X1 U1584 ( .A(\mem<8><4> ), .B(n1262), .Y(n1684) );
  OAI21X1 U1585 ( .A(n1261), .B(n1276), .C(n1684), .Y(n1971) );
  NAND2X1 U1586 ( .A(\mem<8><5> ), .B(n1262), .Y(n1685) );
  OAI21X1 U1587 ( .A(n1261), .B(n1278), .C(n1685), .Y(n1970) );
  NAND2X1 U1588 ( .A(\mem<8><6> ), .B(n1262), .Y(n1686) );
  OAI21X1 U1589 ( .A(n1261), .B(n1279), .C(n1686), .Y(n1969) );
  NAND2X1 U1590 ( .A(\mem<8><7> ), .B(n1262), .Y(n1687) );
  OAI21X1 U1591 ( .A(n1261), .B(n1280), .C(n1687), .Y(n1968) );
  NAND2X1 U1592 ( .A(\mem<8><8> ), .B(n1263), .Y(n1688) );
  OAI21X1 U1593 ( .A(n1261), .B(n1281), .C(n1688), .Y(n1967) );
  NAND2X1 U1594 ( .A(\mem<8><9> ), .B(n1263), .Y(n1689) );
  OAI21X1 U1595 ( .A(n1261), .B(n1283), .C(n1689), .Y(n1966) );
  NAND2X1 U1596 ( .A(\mem<8><10> ), .B(n1263), .Y(n1690) );
  OAI21X1 U1597 ( .A(n1261), .B(n1284), .C(n1690), .Y(n1965) );
  NAND2X1 U1598 ( .A(\mem<8><11> ), .B(n1263), .Y(n1691) );
  OAI21X1 U1599 ( .A(n1261), .B(n1285), .C(n1691), .Y(n1964) );
  NAND2X1 U1600 ( .A(\mem<8><12> ), .B(n1263), .Y(n1692) );
  OAI21X1 U1601 ( .A(n1261), .B(n1287), .C(n1692), .Y(n1963) );
  NAND2X1 U1602 ( .A(\mem<8><13> ), .B(n1263), .Y(n1693) );
  OAI21X1 U1603 ( .A(n1261), .B(n1289), .C(n1693), .Y(n1962) );
  NAND2X1 U1604 ( .A(\mem<8><14> ), .B(n1263), .Y(n1694) );
  OAI21X1 U1605 ( .A(n1261), .B(n1291), .C(n1694), .Y(n1961) );
  NAND2X1 U1606 ( .A(\mem<8><15> ), .B(n1263), .Y(n1695) );
  OAI21X1 U1607 ( .A(n1261), .B(n1293), .C(n1695), .Y(n1960) );
  NAND3X1 U1608 ( .A(n1300), .B(n2344), .C(n1302), .Y(n1696) );
  NAND2X1 U1609 ( .A(\mem<7><0> ), .B(n140), .Y(n1697) );
  OAI21X1 U1610 ( .A(n139), .B(n1271), .C(n1697), .Y(n1959) );
  NAND2X1 U1611 ( .A(\mem<7><1> ), .B(n140), .Y(n1698) );
  OAI21X1 U1612 ( .A(n139), .B(n1273), .C(n1698), .Y(n1958) );
  NAND2X1 U1613 ( .A(\mem<7><2> ), .B(n140), .Y(n1699) );
  OAI21X1 U1614 ( .A(n139), .B(n1274), .C(n1699), .Y(n1957) );
  NAND2X1 U1615 ( .A(\mem<7><3> ), .B(n140), .Y(n1700) );
  OAI21X1 U1616 ( .A(n139), .B(n1275), .C(n1700), .Y(n1956) );
  NAND2X1 U1617 ( .A(\mem<7><4> ), .B(n140), .Y(n1701) );
  OAI21X1 U1618 ( .A(n139), .B(n1276), .C(n1701), .Y(n1955) );
  NAND2X1 U1619 ( .A(\mem<7><5> ), .B(n140), .Y(n1702) );
  OAI21X1 U1620 ( .A(n139), .B(n1278), .C(n1702), .Y(n1954) );
  NAND2X1 U1621 ( .A(\mem<7><6> ), .B(n140), .Y(n1703) );
  OAI21X1 U1622 ( .A(n139), .B(n1279), .C(n1703), .Y(n1953) );
  NAND2X1 U1623 ( .A(\mem<7><7> ), .B(n140), .Y(n1704) );
  OAI21X1 U1624 ( .A(n139), .B(n1280), .C(n1704), .Y(n1952) );
  NAND2X1 U1625 ( .A(\mem<7><8> ), .B(n140), .Y(n1705) );
  OAI21X1 U1626 ( .A(n139), .B(n1281), .C(n1705), .Y(n1951) );
  NAND2X1 U1627 ( .A(\mem<7><9> ), .B(n140), .Y(n1706) );
  OAI21X1 U1628 ( .A(n139), .B(n1283), .C(n1706), .Y(n1950) );
  NAND2X1 U1629 ( .A(\mem<7><10> ), .B(n140), .Y(n1707) );
  OAI21X1 U1630 ( .A(n139), .B(n1284), .C(n1707), .Y(n1949) );
  NAND2X1 U1631 ( .A(\mem<7><11> ), .B(n140), .Y(n1708) );
  OAI21X1 U1632 ( .A(n139), .B(n1285), .C(n1708), .Y(n1948) );
  NAND2X1 U1633 ( .A(\mem<7><12> ), .B(n140), .Y(n1709) );
  OAI21X1 U1634 ( .A(n139), .B(n1287), .C(n1709), .Y(n1947) );
  NAND2X1 U1635 ( .A(\mem<7><13> ), .B(n140), .Y(n1710) );
  OAI21X1 U1636 ( .A(n139), .B(n1289), .C(n1710), .Y(n1946) );
  NAND2X1 U1637 ( .A(\mem<7><14> ), .B(n140), .Y(n1711) );
  OAI21X1 U1638 ( .A(n139), .B(n1291), .C(n1711), .Y(n1945) );
  NAND2X1 U1639 ( .A(\mem<7><15> ), .B(n140), .Y(n1712) );
  OAI21X1 U1640 ( .A(n139), .B(n1293), .C(n1712), .Y(n1944) );
  NAND2X1 U1641 ( .A(\mem<6><0> ), .B(n143), .Y(n1713) );
  OAI21X1 U1642 ( .A(n142), .B(n1272), .C(n1713), .Y(n1943) );
  NAND2X1 U1643 ( .A(\mem<6><1> ), .B(n143), .Y(n1714) );
  OAI21X1 U1644 ( .A(n142), .B(n1273), .C(n1714), .Y(n1942) );
  NAND2X1 U1645 ( .A(\mem<6><2> ), .B(n143), .Y(n1715) );
  OAI21X1 U1646 ( .A(n142), .B(n1274), .C(n1715), .Y(n1941) );
  NAND2X1 U1647 ( .A(\mem<6><3> ), .B(n143), .Y(n1716) );
  OAI21X1 U1648 ( .A(n142), .B(n1275), .C(n1716), .Y(n1940) );
  NAND2X1 U1649 ( .A(\mem<6><4> ), .B(n143), .Y(n1717) );
  OAI21X1 U1650 ( .A(n142), .B(n1276), .C(n1717), .Y(n1939) );
  NAND2X1 U1651 ( .A(\mem<6><5> ), .B(n143), .Y(n1718) );
  OAI21X1 U1652 ( .A(n142), .B(n1278), .C(n1718), .Y(n1938) );
  NAND2X1 U1653 ( .A(\mem<6><6> ), .B(n143), .Y(n1719) );
  OAI21X1 U1654 ( .A(n142), .B(n1279), .C(n1719), .Y(n1937) );
  NAND2X1 U1655 ( .A(\mem<6><7> ), .B(n143), .Y(n1720) );
  OAI21X1 U1656 ( .A(n142), .B(n1280), .C(n1720), .Y(n1936) );
  NAND2X1 U1657 ( .A(\mem<6><8> ), .B(n143), .Y(n1721) );
  OAI21X1 U1658 ( .A(n142), .B(n1281), .C(n1721), .Y(n1935) );
  NAND2X1 U1659 ( .A(\mem<6><9> ), .B(n143), .Y(n1722) );
  OAI21X1 U1660 ( .A(n142), .B(n1283), .C(n1722), .Y(n1934) );
  NAND2X1 U1661 ( .A(\mem<6><10> ), .B(n143), .Y(n1723) );
  OAI21X1 U1662 ( .A(n142), .B(n1284), .C(n1723), .Y(n1933) );
  NAND2X1 U1663 ( .A(\mem<6><11> ), .B(n143), .Y(n1724) );
  OAI21X1 U1664 ( .A(n142), .B(n1285), .C(n1724), .Y(n1932) );
  NAND2X1 U1665 ( .A(\mem<6><12> ), .B(n143), .Y(n1725) );
  OAI21X1 U1666 ( .A(n142), .B(n1287), .C(n1725), .Y(n1931) );
  NAND2X1 U1667 ( .A(\mem<6><13> ), .B(n143), .Y(n1726) );
  OAI21X1 U1668 ( .A(n142), .B(n1289), .C(n1726), .Y(n1930) );
  NAND2X1 U1669 ( .A(\mem<6><14> ), .B(n143), .Y(n1727) );
  OAI21X1 U1670 ( .A(n142), .B(n1291), .C(n1727), .Y(n1929) );
  NAND2X1 U1671 ( .A(\mem<6><15> ), .B(n143), .Y(n1728) );
  OAI21X1 U1672 ( .A(n142), .B(n1293), .C(n1728), .Y(n1928) );
  NAND2X1 U1673 ( .A(\mem<5><0> ), .B(n147), .Y(n1730) );
  OAI21X1 U1674 ( .A(n145), .B(n1271), .C(n1730), .Y(n1927) );
  NAND2X1 U1675 ( .A(\mem<5><1> ), .B(n147), .Y(n1731) );
  OAI21X1 U1676 ( .A(n145), .B(n1273), .C(n1731), .Y(n1926) );
  NAND2X1 U1677 ( .A(\mem<5><2> ), .B(n147), .Y(n1732) );
  OAI21X1 U1678 ( .A(n145), .B(n1274), .C(n1732), .Y(n1925) );
  NAND2X1 U1679 ( .A(\mem<5><3> ), .B(n147), .Y(n1733) );
  OAI21X1 U1680 ( .A(n145), .B(n1275), .C(n1733), .Y(n1924) );
  NAND2X1 U1681 ( .A(\mem<5><4> ), .B(n147), .Y(n1734) );
  OAI21X1 U1682 ( .A(n145), .B(n1276), .C(n1734), .Y(n1923) );
  NAND2X1 U1683 ( .A(\mem<5><5> ), .B(n147), .Y(n1735) );
  OAI21X1 U1684 ( .A(n145), .B(n1278), .C(n1735), .Y(n1922) );
  NAND2X1 U1685 ( .A(\mem<5><6> ), .B(n147), .Y(n1736) );
  OAI21X1 U1686 ( .A(n145), .B(n1279), .C(n1736), .Y(n1921) );
  NAND2X1 U1687 ( .A(\mem<5><7> ), .B(n147), .Y(n1737) );
  OAI21X1 U1688 ( .A(n145), .B(n1280), .C(n1737), .Y(n1920) );
  NAND2X1 U1689 ( .A(\mem<5><8> ), .B(n146), .Y(n1738) );
  OAI21X1 U1690 ( .A(n145), .B(n1281), .C(n1738), .Y(n1919) );
  NAND2X1 U1691 ( .A(\mem<5><9> ), .B(n146), .Y(n1739) );
  OAI21X1 U1692 ( .A(n145), .B(n1283), .C(n1739), .Y(n1918) );
  NAND2X1 U1693 ( .A(\mem<5><10> ), .B(n146), .Y(n1740) );
  OAI21X1 U1694 ( .A(n145), .B(n1284), .C(n1740), .Y(n1917) );
  NAND2X1 U1695 ( .A(\mem<5><11> ), .B(n146), .Y(n1741) );
  OAI21X1 U1696 ( .A(n145), .B(n1285), .C(n1741), .Y(n1916) );
  NAND2X1 U1697 ( .A(\mem<5><12> ), .B(n146), .Y(n1742) );
  OAI21X1 U1698 ( .A(n145), .B(n1287), .C(n1742), .Y(n1915) );
  NAND2X1 U1699 ( .A(\mem<5><13> ), .B(n146), .Y(n1743) );
  OAI21X1 U1700 ( .A(n145), .B(n1289), .C(n1743), .Y(n1914) );
  NAND2X1 U1701 ( .A(\mem<5><14> ), .B(n146), .Y(n1744) );
  OAI21X1 U1702 ( .A(n145), .B(n1291), .C(n1744), .Y(n1913) );
  NAND2X1 U1703 ( .A(\mem<5><15> ), .B(n146), .Y(n1745) );
  OAI21X1 U1704 ( .A(n145), .B(n1293), .C(n1745), .Y(n1912) );
  NAND2X1 U1705 ( .A(\mem<4><0> ), .B(n151), .Y(n1747) );
  OAI21X1 U1706 ( .A(n149), .B(n1272), .C(n1747), .Y(n1911) );
  NAND2X1 U1707 ( .A(\mem<4><1> ), .B(n151), .Y(n1748) );
  OAI21X1 U1708 ( .A(n149), .B(n1273), .C(n1748), .Y(n1910) );
  NAND2X1 U1709 ( .A(\mem<4><2> ), .B(n151), .Y(n1749) );
  OAI21X1 U1710 ( .A(n149), .B(n1274), .C(n1749), .Y(n1909) );
  NAND2X1 U1711 ( .A(\mem<4><3> ), .B(n151), .Y(n1750) );
  OAI21X1 U1712 ( .A(n149), .B(n1275), .C(n1750), .Y(n1908) );
  NAND2X1 U1713 ( .A(\mem<4><4> ), .B(n151), .Y(n1751) );
  OAI21X1 U1714 ( .A(n149), .B(n1276), .C(n1751), .Y(n1907) );
  NAND2X1 U1715 ( .A(\mem<4><5> ), .B(n151), .Y(n1752) );
  OAI21X1 U1716 ( .A(n149), .B(n1278), .C(n1752), .Y(n1906) );
  NAND2X1 U1717 ( .A(\mem<4><6> ), .B(n151), .Y(n1753) );
  OAI21X1 U1718 ( .A(n149), .B(n1279), .C(n1753), .Y(n1905) );
  NAND2X1 U1719 ( .A(\mem<4><7> ), .B(n151), .Y(n1754) );
  OAI21X1 U1720 ( .A(n149), .B(n1280), .C(n1754), .Y(n1904) );
  NAND2X1 U1721 ( .A(\mem<4><8> ), .B(n150), .Y(n1755) );
  OAI21X1 U1722 ( .A(n149), .B(n1281), .C(n1755), .Y(n1903) );
  NAND2X1 U1723 ( .A(\mem<4><9> ), .B(n150), .Y(n1756) );
  OAI21X1 U1724 ( .A(n149), .B(n1283), .C(n1756), .Y(n1902) );
  NAND2X1 U1725 ( .A(\mem<4><10> ), .B(n150), .Y(n1757) );
  OAI21X1 U1726 ( .A(n149), .B(n1284), .C(n1757), .Y(n1901) );
  NAND2X1 U1727 ( .A(\mem<4><11> ), .B(n150), .Y(n1758) );
  OAI21X1 U1728 ( .A(n149), .B(n1285), .C(n1758), .Y(n1900) );
  NAND2X1 U1729 ( .A(\mem<4><12> ), .B(n150), .Y(n1759) );
  OAI21X1 U1730 ( .A(n149), .B(n1287), .C(n1759), .Y(n1899) );
  NAND2X1 U1731 ( .A(\mem<4><13> ), .B(n150), .Y(n1760) );
  OAI21X1 U1732 ( .A(n149), .B(n1289), .C(n1760), .Y(n1898) );
  NAND2X1 U1733 ( .A(\mem<4><14> ), .B(n150), .Y(n1761) );
  OAI21X1 U1734 ( .A(n149), .B(n1291), .C(n1761), .Y(n1897) );
  NAND2X1 U1735 ( .A(\mem<4><15> ), .B(n150), .Y(n1762) );
  OAI21X1 U1736 ( .A(n149), .B(n1293), .C(n1762), .Y(n1896) );
  NAND2X1 U1737 ( .A(\mem<3><0> ), .B(n155), .Y(n1764) );
  OAI21X1 U1738 ( .A(n153), .B(n1271), .C(n1764), .Y(n1895) );
  NAND2X1 U1739 ( .A(\mem<3><1> ), .B(n155), .Y(n1765) );
  OAI21X1 U1740 ( .A(n153), .B(n1273), .C(n1765), .Y(n1894) );
  NAND2X1 U1741 ( .A(\mem<3><2> ), .B(n155), .Y(n1766) );
  OAI21X1 U1742 ( .A(n153), .B(n1274), .C(n1766), .Y(n1893) );
  NAND2X1 U1743 ( .A(\mem<3><3> ), .B(n155), .Y(n1767) );
  OAI21X1 U1744 ( .A(n153), .B(n1275), .C(n1767), .Y(n1892) );
  NAND2X1 U1745 ( .A(\mem<3><4> ), .B(n155), .Y(n1768) );
  OAI21X1 U1746 ( .A(n153), .B(n1276), .C(n1768), .Y(n1891) );
  NAND2X1 U1747 ( .A(\mem<3><5> ), .B(n155), .Y(n1769) );
  OAI21X1 U1748 ( .A(n153), .B(n1278), .C(n1769), .Y(n1890) );
  NAND2X1 U1749 ( .A(\mem<3><6> ), .B(n155), .Y(n1770) );
  OAI21X1 U1750 ( .A(n153), .B(n1279), .C(n1770), .Y(n1889) );
  NAND2X1 U1751 ( .A(\mem<3><7> ), .B(n155), .Y(n1771) );
  OAI21X1 U1752 ( .A(n153), .B(n1280), .C(n1771), .Y(n1888) );
  NAND2X1 U1753 ( .A(\mem<3><8> ), .B(n154), .Y(n1772) );
  OAI21X1 U1754 ( .A(n153), .B(n1281), .C(n1772), .Y(n1887) );
  NAND2X1 U1755 ( .A(\mem<3><9> ), .B(n154), .Y(n1773) );
  OAI21X1 U1756 ( .A(n153), .B(n1283), .C(n1773), .Y(n1886) );
  NAND2X1 U1757 ( .A(\mem<3><10> ), .B(n154), .Y(n1774) );
  OAI21X1 U1758 ( .A(n153), .B(n1284), .C(n1774), .Y(n1885) );
  NAND2X1 U1759 ( .A(\mem<3><11> ), .B(n154), .Y(n1775) );
  OAI21X1 U1760 ( .A(n153), .B(n1285), .C(n1775), .Y(n1884) );
  NAND2X1 U1761 ( .A(\mem<3><12> ), .B(n154), .Y(n1776) );
  OAI21X1 U1762 ( .A(n153), .B(n1287), .C(n1776), .Y(n1883) );
  NAND2X1 U1763 ( .A(\mem<3><13> ), .B(n154), .Y(n1777) );
  OAI21X1 U1764 ( .A(n153), .B(n1289), .C(n1777), .Y(n1882) );
  NAND2X1 U1765 ( .A(\mem<3><14> ), .B(n154), .Y(n1778) );
  OAI21X1 U1766 ( .A(n153), .B(n1291), .C(n1778), .Y(n1881) );
  NAND2X1 U1767 ( .A(\mem<3><15> ), .B(n154), .Y(n1779) );
  OAI21X1 U1768 ( .A(n153), .B(n1293), .C(n1779), .Y(n1880) );
  NAND2X1 U1769 ( .A(\mem<2><0> ), .B(n159), .Y(n1781) );
  OAI21X1 U1770 ( .A(n157), .B(n1272), .C(n1781), .Y(n1879) );
  NAND2X1 U1771 ( .A(\mem<2><1> ), .B(n159), .Y(n1782) );
  OAI21X1 U1772 ( .A(n157), .B(n1273), .C(n1782), .Y(n1878) );
  NAND2X1 U1773 ( .A(\mem<2><2> ), .B(n159), .Y(n1783) );
  OAI21X1 U1774 ( .A(n157), .B(n1274), .C(n1783), .Y(n1877) );
  NAND2X1 U1775 ( .A(\mem<2><3> ), .B(n159), .Y(n1784) );
  OAI21X1 U1776 ( .A(n157), .B(n1275), .C(n1784), .Y(n1876) );
  NAND2X1 U1777 ( .A(\mem<2><4> ), .B(n159), .Y(n1785) );
  OAI21X1 U1778 ( .A(n157), .B(n1276), .C(n1785), .Y(n1875) );
  NAND2X1 U1779 ( .A(\mem<2><5> ), .B(n159), .Y(n1786) );
  OAI21X1 U1780 ( .A(n157), .B(n1278), .C(n1786), .Y(n1874) );
  NAND2X1 U1781 ( .A(\mem<2><6> ), .B(n159), .Y(n1787) );
  OAI21X1 U1782 ( .A(n157), .B(n1279), .C(n1787), .Y(n1873) );
  NAND2X1 U1783 ( .A(\mem<2><7> ), .B(n159), .Y(n1788) );
  OAI21X1 U1784 ( .A(n157), .B(n1280), .C(n1788), .Y(n1872) );
  NAND2X1 U1785 ( .A(\mem<2><8> ), .B(n158), .Y(n1789) );
  OAI21X1 U1786 ( .A(n157), .B(n1281), .C(n1789), .Y(n1871) );
  NAND2X1 U1787 ( .A(\mem<2><9> ), .B(n158), .Y(n1790) );
  OAI21X1 U1788 ( .A(n157), .B(n1283), .C(n1790), .Y(n1870) );
  NAND2X1 U1789 ( .A(\mem<2><10> ), .B(n158), .Y(n1791) );
  OAI21X1 U1790 ( .A(n157), .B(n1284), .C(n1791), .Y(n1869) );
  NAND2X1 U1791 ( .A(\mem<2><11> ), .B(n158), .Y(n1792) );
  OAI21X1 U1792 ( .A(n157), .B(n1285), .C(n1792), .Y(n1868) );
  NAND2X1 U1793 ( .A(\mem<2><12> ), .B(n158), .Y(n1793) );
  OAI21X1 U1794 ( .A(n157), .B(n1287), .C(n1793), .Y(n1867) );
  NAND2X1 U1795 ( .A(\mem<2><13> ), .B(n158), .Y(n1794) );
  OAI21X1 U1796 ( .A(n157), .B(n1289), .C(n1794), .Y(n1866) );
  NAND2X1 U1797 ( .A(\mem<2><14> ), .B(n158), .Y(n1795) );
  OAI21X1 U1798 ( .A(n157), .B(n1291), .C(n1795), .Y(n1865) );
  NAND2X1 U1799 ( .A(\mem<2><15> ), .B(n158), .Y(n1796) );
  OAI21X1 U1800 ( .A(n157), .B(n1293), .C(n1796), .Y(n1864) );
  NAND2X1 U1801 ( .A(\mem<1><0> ), .B(n163), .Y(n1798) );
  OAI21X1 U1802 ( .A(n161), .B(n1271), .C(n1798), .Y(n1863) );
  NAND2X1 U1803 ( .A(\mem<1><1> ), .B(n163), .Y(n1799) );
  OAI21X1 U1804 ( .A(n161), .B(n1273), .C(n1799), .Y(n1862) );
  NAND2X1 U1805 ( .A(\mem<1><2> ), .B(n163), .Y(n1800) );
  OAI21X1 U1806 ( .A(n161), .B(n1274), .C(n1800), .Y(n1861) );
  NAND2X1 U1807 ( .A(\mem<1><3> ), .B(n163), .Y(n1801) );
  OAI21X1 U1808 ( .A(n161), .B(n1275), .C(n1801), .Y(n1860) );
  NAND2X1 U1809 ( .A(\mem<1><4> ), .B(n163), .Y(n1802) );
  OAI21X1 U1810 ( .A(n161), .B(n1276), .C(n1802), .Y(n1859) );
  NAND2X1 U1811 ( .A(\mem<1><5> ), .B(n163), .Y(n1803) );
  OAI21X1 U1812 ( .A(n161), .B(n1278), .C(n1803), .Y(n1858) );
  NAND2X1 U1813 ( .A(\mem<1><6> ), .B(n163), .Y(n1804) );
  OAI21X1 U1814 ( .A(n161), .B(n1279), .C(n1804), .Y(n1857) );
  NAND2X1 U1815 ( .A(\mem<1><7> ), .B(n163), .Y(n1805) );
  OAI21X1 U1816 ( .A(n161), .B(n1280), .C(n1805), .Y(n1856) );
  NAND2X1 U1817 ( .A(\mem<1><8> ), .B(n162), .Y(n1806) );
  OAI21X1 U1818 ( .A(n161), .B(n1281), .C(n1806), .Y(n1855) );
  NAND2X1 U1819 ( .A(\mem<1><9> ), .B(n162), .Y(n1807) );
  OAI21X1 U1820 ( .A(n161), .B(n1283), .C(n1807), .Y(n1854) );
  NAND2X1 U1821 ( .A(\mem<1><10> ), .B(n162), .Y(n1808) );
  OAI21X1 U1822 ( .A(n161), .B(n1284), .C(n1808), .Y(n1853) );
  NAND2X1 U1823 ( .A(\mem<1><11> ), .B(n162), .Y(n1809) );
  OAI21X1 U1824 ( .A(n161), .B(n1285), .C(n1809), .Y(n1852) );
  NAND2X1 U1825 ( .A(\mem<1><12> ), .B(n162), .Y(n1810) );
  OAI21X1 U1826 ( .A(n161), .B(n1287), .C(n1810), .Y(n1851) );
  NAND2X1 U1827 ( .A(\mem<1><13> ), .B(n162), .Y(n1811) );
  OAI21X1 U1828 ( .A(n161), .B(n1289), .C(n1811), .Y(n1850) );
  NAND2X1 U1829 ( .A(\mem<1><14> ), .B(n162), .Y(n1812) );
  OAI21X1 U1830 ( .A(n161), .B(n1291), .C(n1812), .Y(n1849) );
  NAND2X1 U1831 ( .A(\mem<1><15> ), .B(n162), .Y(n1813) );
  OAI21X1 U1832 ( .A(n161), .B(n1293), .C(n1813), .Y(n1848) );
  NAND2X1 U1833 ( .A(\mem<0><0> ), .B(n1265), .Y(n1816) );
  OAI21X1 U1834 ( .A(n1264), .B(n1272), .C(n1816), .Y(n1847) );
  NAND2X1 U1835 ( .A(\mem<0><1> ), .B(n1265), .Y(n1817) );
  OAI21X1 U1836 ( .A(n1264), .B(n1273), .C(n1817), .Y(n1846) );
  NAND2X1 U1837 ( .A(\mem<0><2> ), .B(n1265), .Y(n1818) );
  OAI21X1 U1838 ( .A(n1264), .B(n1274), .C(n1818), .Y(n1845) );
  NAND2X1 U1839 ( .A(\mem<0><3> ), .B(n1265), .Y(n1819) );
  OAI21X1 U1840 ( .A(n1264), .B(n1275), .C(n1819), .Y(n1844) );
  NAND2X1 U1841 ( .A(\mem<0><4> ), .B(n1265), .Y(n1820) );
  OAI21X1 U1842 ( .A(n1264), .B(n1276), .C(n1820), .Y(n1843) );
  NAND2X1 U1843 ( .A(\mem<0><5> ), .B(n1265), .Y(n1821) );
  OAI21X1 U1844 ( .A(n1264), .B(n1278), .C(n1821), .Y(n1842) );
  NAND2X1 U1845 ( .A(\mem<0><6> ), .B(n1265), .Y(n1822) );
  OAI21X1 U1846 ( .A(n1264), .B(n1279), .C(n1822), .Y(n1841) );
  NAND2X1 U1847 ( .A(\mem<0><7> ), .B(n1265), .Y(n1823) );
  OAI21X1 U1848 ( .A(n1264), .B(n1280), .C(n1823), .Y(n1840) );
  NAND2X1 U1849 ( .A(\mem<0><8> ), .B(n1266), .Y(n1824) );
  OAI21X1 U1850 ( .A(n1264), .B(n1281), .C(n1824), .Y(n1839) );
  NAND2X1 U1851 ( .A(\mem<0><9> ), .B(n1266), .Y(n1825) );
  OAI21X1 U1852 ( .A(n1264), .B(n1283), .C(n1825), .Y(n1838) );
  NAND2X1 U1853 ( .A(\mem<0><10> ), .B(n1266), .Y(n1826) );
  OAI21X1 U1854 ( .A(n1264), .B(n1284), .C(n1826), .Y(n1837) );
  NAND2X1 U1855 ( .A(\mem<0><11> ), .B(n1266), .Y(n1827) );
  OAI21X1 U1856 ( .A(n1264), .B(n1285), .C(n1827), .Y(n1836) );
  NAND2X1 U1857 ( .A(\mem<0><12> ), .B(n1266), .Y(n1828) );
  OAI21X1 U1858 ( .A(n1264), .B(n1287), .C(n1828), .Y(n1835) );
  NAND2X1 U1859 ( .A(\mem<0><13> ), .B(n1266), .Y(n1829) );
  OAI21X1 U1860 ( .A(n1264), .B(n1289), .C(n1829), .Y(n1834) );
  NAND2X1 U1861 ( .A(\mem<0><14> ), .B(n1266), .Y(n1830) );
  OAI21X1 U1862 ( .A(n1264), .B(n1291), .C(n1830), .Y(n1833) );
  NAND2X1 U1863 ( .A(\mem<0><15> ), .B(n1266), .Y(n1831) );
  OAI21X1 U1864 ( .A(n1264), .B(n1293), .C(n1831), .Y(n1832) );
endmodule


module memc_Size5 ( .data_out({\data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        write, clk, rst, createdump, .file_id({\file_id<4> , \file_id<3> , 
        \file_id<2> , \file_id<1> , \file_id<0> }) );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<4> , \data_in<3> , \data_in<2> ,
         \data_in<1> , \data_in<0> , write, clk, rst, createdump, \file_id<4> ,
         \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> ;
  output \data_out<4> , \data_out<3> , \data_out<2> , \data_out<1> ,
         \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><4> , \mem<0><3> , \mem<0><2> ,
         \mem<0><1> , \mem<0><0> , \mem<1><4> , \mem<1><3> , \mem<1><2> ,
         \mem<1><1> , \mem<1><0> , \mem<2><4> , \mem<2><3> , \mem<2><2> ,
         \mem<2><1> , \mem<2><0> , \mem<3><4> , \mem<3><3> , \mem<3><2> ,
         \mem<3><1> , \mem<3><0> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><4> , \mem<5><3> , \mem<5><2> ,
         \mem<5><1> , \mem<5><0> , \mem<6><4> , \mem<6><3> , \mem<6><2> ,
         \mem<6><1> , \mem<6><0> , \mem<7><4> , \mem<7><3> , \mem<7><2> ,
         \mem<7><1> , \mem<7><0> , \mem<8><4> , \mem<8><3> , \mem<8><2> ,
         \mem<8><1> , \mem<8><0> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><4> , \mem<10><3> , \mem<10><2> ,
         \mem<10><1> , \mem<10><0> , \mem<11><4> , \mem<11><3> , \mem<11><2> ,
         \mem<11><1> , \mem<11><0> , \mem<12><4> , \mem<12><3> , \mem<12><2> ,
         \mem<12><1> , \mem<12><0> , \mem<13><4> , \mem<13><3> , \mem<13><2> ,
         \mem<13><1> , \mem<13><0> , \mem<14><4> , \mem<14><3> , \mem<14><2> ,
         \mem<14><1> , \mem<14><0> , \mem<15><4> , \mem<15><3> , \mem<15><2> ,
         \mem<15><1> , \mem<15><0> , \mem<16><4> , \mem<16><3> , \mem<16><2> ,
         \mem<16><1> , \mem<16><0> , \mem<17><4> , \mem<17><3> , \mem<17><2> ,
         \mem<17><1> , \mem<17><0> , \mem<18><4> , \mem<18><3> , \mem<18><2> ,
         \mem<18><1> , \mem<18><0> , \mem<19><4> , \mem<19><3> , \mem<19><2> ,
         \mem<19><1> , \mem<19><0> , \mem<20><4> , \mem<20><3> , \mem<20><2> ,
         \mem<20><1> , \mem<20><0> , \mem<21><4> , \mem<21><3> , \mem<21><2> ,
         \mem<21><1> , \mem<21><0> , \mem<22><4> , \mem<22><3> , \mem<22><2> ,
         \mem<22><1> , \mem<22><0> , \mem<23><4> , \mem<23><3> , \mem<23><2> ,
         \mem<23><1> , \mem<23><0> , \mem<24><4> , \mem<24><3> , \mem<24><2> ,
         \mem<24><1> , \mem<24><0> , \mem<25><4> , \mem<25><3> , \mem<25><2> ,
         \mem<25><1> , \mem<25><0> , \mem<26><4> , \mem<26><3> , \mem<26><2> ,
         \mem<26><1> , \mem<26><0> , \mem<27><4> , \mem<27><3> , \mem<27><2> ,
         \mem<27><1> , \mem<27><0> , \mem<28><4> , \mem<28><3> , \mem<28><2> ,
         \mem<28><1> , \mem<28><0> , \mem<29><4> , \mem<29><3> , \mem<29><2> ,
         \mem<29><1> , \mem<29><0> , \mem<30><4> , \mem<30><3> , \mem<30><2> ,
         \mem<30><1> , \mem<30><0> , \mem<31><4> , \mem<31><3> , \mem<31><2> ,
         \mem<31><1> , \mem<31><0> , N17, N18, N19, N20, N21, n56, n57, n65,
         n73, n81, n89, n97, n105, n113, n114, n115, n136, n172, n229, n286,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n58, n59, n60, n61, n62, n63, n64, n66, n67,
         n68, n69, n70, n71, n72, n74, n75, n76, n77, n78, n79, n80, n82, n83,
         n84, n85, n86, n87, n88, n90, n91, n92, n93, n94, n95, n96, n98, n99,
         n100, n101, n102, n103, n104, n106, n107, n108, n109, n110, n111,
         n112, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n287, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><4>  ( .D(n447), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n446), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n445), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n444), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n443), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n442), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n441), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n440), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n439), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n438), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n437), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n436), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n435), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n434), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n433), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n432), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n431), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n430), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n429), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n428), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n427), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n426), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n425), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n424), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n423), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n422), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n421), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n420), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n419), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n418), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n417), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n416), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n415), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n414), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n413), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n412), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n411), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n410), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n409), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n408), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n407), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n406), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n405), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n404), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n403), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n402), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n401), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n400), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n399), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n398), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n397), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n396), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n395), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n394), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n393), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n392), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n391), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n390), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n389), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n388), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n387), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n386), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n385), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n384), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n383), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n382), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n381), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n380), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n379), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n378), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n377), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n376), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n375), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n374), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n373), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n372), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n371), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n370), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n369), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n368), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n367), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n366), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n365), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n364), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n363), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n362), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n361), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n360), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n359), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n358), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n357), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n356), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n355), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n354), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n353), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n352), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n351), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n350), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n349), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n348), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n347), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n346), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n345), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n344), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n343), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n342), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n341), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n340), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n339), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n338), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n337), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n336), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n335), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n334), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n333), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n332), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n331), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n330), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n329), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n328), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n327), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n326), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n325), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n324), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n323), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n322), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n321), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n320), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n319), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n318), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n317), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n316), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n315), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n314), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n313), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n312), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n311), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n310), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n309), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n308), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n307), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n306), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n305), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n304), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n303), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n302), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n301), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n300), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n299), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n298), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n297), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n296), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n295), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n294), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n293), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n292), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n291), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n290), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n289), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n288), .CLK(clk), .Q(\mem<31><0> ) );
  AND2X2 U2 ( .A(write), .B(n816), .Y(n56) );
  OAI21X1 U50 ( .A(n571), .B(n815), .C(n496), .Y(n288) );
  OAI21X1 U52 ( .A(n571), .B(n814), .C(n494), .Y(n289) );
  OAI21X1 U54 ( .A(n571), .B(n813), .C(n492), .Y(n290) );
  OAI21X1 U56 ( .A(n571), .B(n812), .C(n490), .Y(n291) );
  OAI21X1 U58 ( .A(n571), .B(n811), .C(n488), .Y(n292) );
  OAI21X1 U62 ( .A(n815), .B(n633), .C(n486), .Y(n293) );
  OAI21X1 U64 ( .A(n814), .B(n633), .C(n484), .Y(n294) );
  OAI21X1 U66 ( .A(n813), .B(n633), .C(n482), .Y(n295) );
  OAI21X1 U68 ( .A(n812), .B(n633), .C(n480), .Y(n296) );
  OAI21X1 U70 ( .A(n811), .B(n633), .C(n478), .Y(n297) );
  OAI21X1 U74 ( .A(n815), .B(n631), .C(n476), .Y(n298) );
  OAI21X1 U76 ( .A(n814), .B(n631), .C(n474), .Y(n299) );
  OAI21X1 U78 ( .A(n813), .B(n631), .C(n472), .Y(n300) );
  OAI21X1 U80 ( .A(n812), .B(n631), .C(n470), .Y(n301) );
  OAI21X1 U82 ( .A(n811), .B(n631), .C(n468), .Y(n302) );
  OAI21X1 U86 ( .A(n815), .B(n629), .C(n466), .Y(n303) );
  OAI21X1 U88 ( .A(n814), .B(n629), .C(n464), .Y(n304) );
  OAI21X1 U90 ( .A(n813), .B(n629), .C(n462), .Y(n305) );
  OAI21X1 U92 ( .A(n812), .B(n629), .C(n460), .Y(n306) );
  OAI21X1 U94 ( .A(n811), .B(n629), .C(n458), .Y(n307) );
  OAI21X1 U98 ( .A(n815), .B(n627), .C(n456), .Y(n308) );
  OAI21X1 U100 ( .A(n814), .B(n627), .C(n454), .Y(n309) );
  OAI21X1 U102 ( .A(n813), .B(n627), .C(n452), .Y(n310) );
  OAI21X1 U104 ( .A(n812), .B(n627), .C(n450), .Y(n311) );
  OAI21X1 U106 ( .A(n811), .B(n627), .C(n448), .Y(n312) );
  OAI21X1 U110 ( .A(n815), .B(n625), .C(n285), .Y(n313) );
  OAI21X1 U112 ( .A(n814), .B(n625), .C(n283), .Y(n314) );
  OAI21X1 U114 ( .A(n813), .B(n625), .C(n281), .Y(n315) );
  OAI21X1 U116 ( .A(n812), .B(n625), .C(n279), .Y(n316) );
  OAI21X1 U118 ( .A(n811), .B(n625), .C(n277), .Y(n317) );
  OAI21X1 U122 ( .A(n815), .B(n623), .C(n275), .Y(n318) );
  OAI21X1 U124 ( .A(n814), .B(n623), .C(n273), .Y(n319) );
  OAI21X1 U126 ( .A(n813), .B(n623), .C(n271), .Y(n320) );
  OAI21X1 U128 ( .A(n812), .B(n623), .C(n269), .Y(n321) );
  OAI21X1 U130 ( .A(n811), .B(n623), .C(n267), .Y(n322) );
  OAI21X1 U134 ( .A(n815), .B(n621), .C(n265), .Y(n323) );
  OAI21X1 U136 ( .A(n814), .B(n621), .C(n263), .Y(n324) );
  OAI21X1 U138 ( .A(n813), .B(n621), .C(n261), .Y(n325) );
  OAI21X1 U140 ( .A(n812), .B(n621), .C(n259), .Y(n326) );
  OAI21X1 U142 ( .A(n811), .B(n621), .C(n257), .Y(n327) );
  NAND3X1 U146 ( .A(N13), .B(n115), .C(N14), .Y(n114) );
  OAI21X1 U147 ( .A(n815), .B(n619), .C(n255), .Y(n328) );
  OAI21X1 U149 ( .A(n814), .B(n619), .C(n253), .Y(n329) );
  OAI21X1 U151 ( .A(n813), .B(n619), .C(n251), .Y(n330) );
  OAI21X1 U153 ( .A(n812), .B(n619), .C(n249), .Y(n331) );
  OAI21X1 U155 ( .A(n811), .B(n619), .C(n247), .Y(n332) );
  OAI21X1 U159 ( .A(n815), .B(n617), .C(n245), .Y(n333) );
  OAI21X1 U161 ( .A(n814), .B(n617), .C(n243), .Y(n334) );
  OAI21X1 U163 ( .A(n813), .B(n617), .C(n241), .Y(n335) );
  OAI21X1 U165 ( .A(n812), .B(n617), .C(n239), .Y(n336) );
  OAI21X1 U167 ( .A(n811), .B(n617), .C(n237), .Y(n337) );
  OAI21X1 U171 ( .A(n815), .B(n615), .C(n235), .Y(n338) );
  OAI21X1 U173 ( .A(n814), .B(n615), .C(n233), .Y(n339) );
  OAI21X1 U175 ( .A(n813), .B(n615), .C(n231), .Y(n340) );
  OAI21X1 U177 ( .A(n812), .B(n615), .C(n228), .Y(n341) );
  OAI21X1 U179 ( .A(n811), .B(n615), .C(n136), .Y(n342) );
  NAND2X1 U180 ( .A(\mem<21><4> ), .B(n549), .Y(n136) );
  OAI21X1 U183 ( .A(n815), .B(n613), .C(n226), .Y(n343) );
  OAI21X1 U185 ( .A(n814), .B(n613), .C(n224), .Y(n344) );
  OAI21X1 U187 ( .A(n813), .B(n613), .C(n222), .Y(n345) );
  OAI21X1 U189 ( .A(n812), .B(n613), .C(n220), .Y(n346) );
  OAI21X1 U191 ( .A(n811), .B(n613), .C(n218), .Y(n347) );
  OAI21X1 U195 ( .A(n815), .B(n611), .C(n216), .Y(n348) );
  OAI21X1 U197 ( .A(n814), .B(n611), .C(n214), .Y(n349) );
  OAI21X1 U199 ( .A(n813), .B(n611), .C(n212), .Y(n350) );
  OAI21X1 U201 ( .A(n812), .B(n611), .C(n210), .Y(n351) );
  OAI21X1 U203 ( .A(n811), .B(n611), .C(n208), .Y(n352) );
  OAI21X1 U207 ( .A(n815), .B(n609), .C(n206), .Y(n353) );
  OAI21X1 U209 ( .A(n814), .B(n609), .C(n204), .Y(n354) );
  OAI21X1 U211 ( .A(n813), .B(n609), .C(n202), .Y(n355) );
  OAI21X1 U213 ( .A(n812), .B(n609), .C(n200), .Y(n356) );
  OAI21X1 U215 ( .A(n811), .B(n609), .C(n198), .Y(n357) );
  OAI21X1 U219 ( .A(n815), .B(n607), .C(n196), .Y(n358) );
  OAI21X1 U221 ( .A(n814), .B(n607), .C(n194), .Y(n359) );
  OAI21X1 U223 ( .A(n813), .B(n607), .C(n192), .Y(n360) );
  OAI21X1 U225 ( .A(n812), .B(n607), .C(n190), .Y(n361) );
  OAI21X1 U227 ( .A(n811), .B(n607), .C(n188), .Y(n362) );
  OAI21X1 U231 ( .A(n815), .B(n605), .C(n186), .Y(n363) );
  OAI21X1 U233 ( .A(n814), .B(n605), .C(n184), .Y(n364) );
  OAI21X1 U235 ( .A(n813), .B(n605), .C(n182), .Y(n365) );
  OAI21X1 U237 ( .A(n812), .B(n605), .C(n180), .Y(n366) );
  OAI21X1 U239 ( .A(n811), .B(n605), .C(n178), .Y(n367) );
  NAND3X1 U243 ( .A(n115), .B(n819), .C(N14), .Y(n172) );
  OAI21X1 U244 ( .A(n815), .B(n603), .C(n176), .Y(n368) );
  OAI21X1 U246 ( .A(n814), .B(n603), .C(n174), .Y(n369) );
  OAI21X1 U248 ( .A(n813), .B(n603), .C(n171), .Y(n370) );
  OAI21X1 U250 ( .A(n812), .B(n603), .C(n169), .Y(n371) );
  OAI21X1 U252 ( .A(n811), .B(n603), .C(n167), .Y(n372) );
  OAI21X1 U256 ( .A(n815), .B(n601), .C(n165), .Y(n373) );
  OAI21X1 U258 ( .A(n814), .B(n601), .C(n163), .Y(n374) );
  OAI21X1 U260 ( .A(n813), .B(n601), .C(n161), .Y(n375) );
  OAI21X1 U262 ( .A(n812), .B(n601), .C(n159), .Y(n376) );
  OAI21X1 U264 ( .A(n811), .B(n601), .C(n157), .Y(n377) );
  OAI21X1 U268 ( .A(n815), .B(n599), .C(n155), .Y(n378) );
  OAI21X1 U270 ( .A(n814), .B(n599), .C(n153), .Y(n379) );
  OAI21X1 U272 ( .A(n813), .B(n599), .C(n151), .Y(n380) );
  OAI21X1 U274 ( .A(n812), .B(n599), .C(n149), .Y(n381) );
  OAI21X1 U276 ( .A(n811), .B(n599), .C(n147), .Y(n382) );
  OAI21X1 U280 ( .A(n815), .B(n597), .C(n145), .Y(n383) );
  OAI21X1 U282 ( .A(n814), .B(n597), .C(n143), .Y(n384) );
  OAI21X1 U284 ( .A(n813), .B(n597), .C(n141), .Y(n385) );
  OAI21X1 U286 ( .A(n812), .B(n597), .C(n139), .Y(n386) );
  OAI21X1 U288 ( .A(n811), .B(n597), .C(n137), .Y(n387) );
  OAI21X1 U292 ( .A(n815), .B(n595), .C(n134), .Y(n388) );
  OAI21X1 U294 ( .A(n814), .B(n595), .C(n132), .Y(n389) );
  OAI21X1 U296 ( .A(n813), .B(n595), .C(n130), .Y(n390) );
  OAI21X1 U298 ( .A(n812), .B(n595), .C(n128), .Y(n391) );
  OAI21X1 U300 ( .A(n811), .B(n595), .C(n126), .Y(n392) );
  OAI21X1 U304 ( .A(n815), .B(n593), .C(n124), .Y(n393) );
  OAI21X1 U306 ( .A(n814), .B(n593), .C(n122), .Y(n394) );
  OAI21X1 U308 ( .A(n813), .B(n593), .C(n120), .Y(n395) );
  OAI21X1 U310 ( .A(n812), .B(n593), .C(n118), .Y(n396) );
  OAI21X1 U312 ( .A(n811), .B(n593), .C(n116), .Y(n397) );
  OAI21X1 U316 ( .A(n815), .B(n591), .C(n111), .Y(n398) );
  OAI21X1 U318 ( .A(n814), .B(n591), .C(n109), .Y(n399) );
  OAI21X1 U320 ( .A(n813), .B(n591), .C(n107), .Y(n400) );
  OAI21X1 U322 ( .A(n812), .B(n591), .C(n104), .Y(n401) );
  OAI21X1 U324 ( .A(n811), .B(n591), .C(n102), .Y(n402) );
  OAI21X1 U328 ( .A(n815), .B(n589), .C(n100), .Y(n403) );
  OAI21X1 U330 ( .A(n814), .B(n589), .C(n98), .Y(n404) );
  OAI21X1 U332 ( .A(n813), .B(n589), .C(n95), .Y(n405) );
  OAI21X1 U334 ( .A(n812), .B(n589), .C(n93), .Y(n406) );
  OAI21X1 U336 ( .A(n811), .B(n589), .C(n91), .Y(n407) );
  NAND3X1 U340 ( .A(n115), .B(n820), .C(N13), .Y(n229) );
  OAI21X1 U341 ( .A(n815), .B(n587), .C(n88), .Y(n408) );
  OAI21X1 U343 ( .A(n814), .B(n587), .C(n86), .Y(n409) );
  OAI21X1 U345 ( .A(n813), .B(n587), .C(n84), .Y(n410) );
  OAI21X1 U347 ( .A(n812), .B(n587), .C(n82), .Y(n411) );
  OAI21X1 U349 ( .A(n811), .B(n587), .C(n79), .Y(n412) );
  NOR3X1 U353 ( .A(n793), .B(n817), .C(n818), .Y(n57) );
  OAI21X1 U354 ( .A(n815), .B(n585), .C(n77), .Y(n413) );
  OAI21X1 U356 ( .A(n814), .B(n585), .C(n75), .Y(n414) );
  OAI21X1 U358 ( .A(n813), .B(n585), .C(n72), .Y(n415) );
  OAI21X1 U360 ( .A(n812), .B(n585), .C(n70), .Y(n416) );
  OAI21X1 U362 ( .A(n811), .B(n585), .C(n68), .Y(n417) );
  NOR3X1 U366 ( .A(n793), .B(n803), .C(n818), .Y(n65) );
  OAI21X1 U367 ( .A(n815), .B(n583), .C(n66), .Y(n418) );
  OAI21X1 U369 ( .A(n814), .B(n583), .C(n63), .Y(n419) );
  OAI21X1 U371 ( .A(n813), .B(n583), .C(n61), .Y(n420) );
  OAI21X1 U373 ( .A(n812), .B(n583), .C(n59), .Y(n421) );
  OAI21X1 U375 ( .A(n811), .B(n583), .C(n55), .Y(n422) );
  NOR3X1 U379 ( .A(n817), .B(n797), .C(n818), .Y(n73) );
  OAI21X1 U380 ( .A(n815), .B(n581), .C(n53), .Y(n423) );
  OAI21X1 U382 ( .A(n814), .B(n581), .C(n51), .Y(n424) );
  OAI21X1 U384 ( .A(n813), .B(n581), .C(n49), .Y(n425) );
  OAI21X1 U386 ( .A(n812), .B(n581), .C(n47), .Y(n426) );
  OAI21X1 U388 ( .A(n811), .B(n581), .C(n45), .Y(n427) );
  NOR3X1 U392 ( .A(n809), .B(n797), .C(n818), .Y(n81) );
  OAI21X1 U393 ( .A(n815), .B(n579), .C(n43), .Y(n428) );
  OAI21X1 U395 ( .A(n814), .B(n579), .C(n41), .Y(n429) );
  OAI21X1 U397 ( .A(n813), .B(n579), .C(n39), .Y(n430) );
  OAI21X1 U399 ( .A(n812), .B(n579), .C(n37), .Y(n431) );
  OAI21X1 U401 ( .A(n811), .B(n579), .C(n35), .Y(n432) );
  NOR3X1 U405 ( .A(n817), .B(N12), .C(n793), .Y(n89) );
  OAI21X1 U406 ( .A(n815), .B(n577), .C(n33), .Y(n433) );
  OAI21X1 U408 ( .A(n814), .B(n577), .C(n31), .Y(n434) );
  OAI21X1 U410 ( .A(n813), .B(n577), .C(n29), .Y(n435) );
  OAI21X1 U412 ( .A(n812), .B(n577), .C(n27), .Y(n436) );
  OAI21X1 U414 ( .A(n811), .B(n577), .C(n25), .Y(n437) );
  NOR3X1 U418 ( .A(n802), .B(N12), .C(n793), .Y(n97) );
  OAI21X1 U419 ( .A(n815), .B(n575), .C(n23), .Y(n438) );
  OAI21X1 U421 ( .A(n814), .B(n575), .C(n21), .Y(n439) );
  OAI21X1 U423 ( .A(n813), .B(n575), .C(n19), .Y(n440) );
  OAI21X1 U425 ( .A(n812), .B(n575), .C(n17), .Y(n441) );
  OAI21X1 U427 ( .A(n811), .B(n575), .C(n15), .Y(n442) );
  NOR3X1 U431 ( .A(n797), .B(N12), .C(n817), .Y(n105) );
  OAI21X1 U432 ( .A(n815), .B(n573), .C(n13), .Y(n443) );
  OAI21X1 U435 ( .A(n814), .B(n573), .C(n11), .Y(n444) );
  OAI21X1 U438 ( .A(n813), .B(n573), .C(n9), .Y(n445) );
  OAI21X1 U441 ( .A(n812), .B(n573), .C(n7), .Y(n446) );
  OAI21X1 U444 ( .A(n811), .B(n573), .C(n5), .Y(n447) );
  NOR3X1 U448 ( .A(n797), .B(N12), .C(n3), .Y(n113) );
  NAND3X1 U449 ( .A(n819), .B(n820), .C(n115), .Y(n286) );
  NOR3X1 U450 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n115) );
  INVX1 U3 ( .A(n788), .Y(N17) );
  AND2X1 U4 ( .A(\mem<31><1> ), .B(n569), .Y(n493) );
  AND2X1 U5 ( .A(\mem<31><2> ), .B(n569), .Y(n491) );
  AND2X1 U6 ( .A(\mem<31><3> ), .B(n569), .Y(n489) );
  AND2X1 U7 ( .A(\mem<31><4> ), .B(n569), .Y(n487) );
  AND2X1 U8 ( .A(\mem<30><2> ), .B(n567), .Y(n481) );
  AND2X1 U9 ( .A(\mem<30><4> ), .B(n567), .Y(n477) );
  AND2X1 U10 ( .A(\mem<29><1> ), .B(n565), .Y(n473) );
  AND2X1 U11 ( .A(\mem<29><2> ), .B(n565), .Y(n471) );
  AND2X1 U12 ( .A(\mem<29><3> ), .B(n565), .Y(n469) );
  AND2X1 U13 ( .A(\mem<29><4> ), .B(n565), .Y(n467) );
  AND2X1 U14 ( .A(\mem<28><2> ), .B(n563), .Y(n461) );
  AND2X1 U15 ( .A(\mem<28><4> ), .B(n563), .Y(n457) );
  AND2X1 U16 ( .A(\mem<27><2> ), .B(n561), .Y(n451) );
  AND2X1 U17 ( .A(\mem<27><4> ), .B(n561), .Y(n287) );
  AND2X1 U18 ( .A(\mem<26><4> ), .B(n559), .Y(n276) );
  AND2X1 U19 ( .A(\mem<25><2> ), .B(n557), .Y(n270) );
  AND2X1 U20 ( .A(\mem<25><4> ), .B(n557), .Y(n266) );
  AND2X1 U21 ( .A(\mem<24><4> ), .B(n555), .Y(n256) );
  AND2X1 U22 ( .A(\mem<23><1> ), .B(n553), .Y(n252) );
  AND2X1 U23 ( .A(\mem<23><2> ), .B(n553), .Y(n250) );
  AND2X1 U24 ( .A(\mem<23><3> ), .B(n553), .Y(n248) );
  AND2X1 U25 ( .A(\mem<23><4> ), .B(n553), .Y(n246) );
  AND2X1 U26 ( .A(\mem<22><2> ), .B(n551), .Y(n240) );
  AND2X1 U27 ( .A(\mem<22><4> ), .B(n551), .Y(n236) );
  AND2X1 U28 ( .A(\mem<21><1> ), .B(n549), .Y(n232) );
  AND2X1 U29 ( .A(\mem<21><2> ), .B(n549), .Y(n230) );
  AND2X1 U30 ( .A(\mem<21><3> ), .B(n549), .Y(n227) );
  AND2X1 U31 ( .A(\mem<20><2> ), .B(n547), .Y(n221) );
  AND2X1 U32 ( .A(\mem<20><4> ), .B(n547), .Y(n217) );
  AND2X1 U33 ( .A(\mem<19><2> ), .B(n545), .Y(n211) );
  AND2X1 U34 ( .A(\mem<19><4> ), .B(n545), .Y(n207) );
  AND2X1 U35 ( .A(\mem<18><4> ), .B(n543), .Y(n197) );
  AND2X1 U36 ( .A(\mem<17><2> ), .B(n541), .Y(n191) );
  AND2X1 U37 ( .A(\mem<17><4> ), .B(n541), .Y(n187) );
  AND2X1 U38 ( .A(\mem<16><4> ), .B(n539), .Y(n177) );
  AND2X1 U39 ( .A(\mem<15><2> ), .B(n537), .Y(n170) );
  AND2X1 U40 ( .A(\mem<15><4> ), .B(n537), .Y(n166) );
  AND2X1 U41 ( .A(\mem<14><4> ), .B(n535), .Y(n156) );
  AND2X1 U42 ( .A(\mem<13><2> ), .B(n533), .Y(n150) );
  AND2X1 U43 ( .A(\mem<13><4> ), .B(n533), .Y(n146) );
  AND2X1 U44 ( .A(\mem<12><4> ), .B(n531), .Y(n135) );
  AND2X1 U45 ( .A(\mem<11><4> ), .B(n529), .Y(n125) );
  AND2X1 U46 ( .A(\mem<10><4> ), .B(n527), .Y(n112) );
  AND2X1 U47 ( .A(\mem<9><4> ), .B(n525), .Y(n101) );
  AND2X1 U48 ( .A(\mem<8><4> ), .B(n523), .Y(n90) );
  AND2X1 U49 ( .A(\mem<7><2> ), .B(n521), .Y(n83) );
  AND2X1 U51 ( .A(\mem<7><4> ), .B(n521), .Y(n78) );
  AND2X1 U53 ( .A(\mem<6><4> ), .B(n519), .Y(n67) );
  AND2X1 U55 ( .A(\mem<5><2> ), .B(n517), .Y(n60) );
  AND2X1 U57 ( .A(\mem<5><4> ), .B(n517), .Y(n54) );
  AND2X1 U59 ( .A(\mem<4><4> ), .B(n515), .Y(n44) );
  AND2X1 U60 ( .A(\mem<3><4> ), .B(n513), .Y(n34) );
  AND2X1 U61 ( .A(\mem<2><4> ), .B(n511), .Y(n24) );
  AND2X1 U63 ( .A(\mem<1><4> ), .B(n509), .Y(n14) );
  AND2X1 U65 ( .A(\mem<0><4> ), .B(n507), .Y(n4) );
  INVX4 U67 ( .A(N11), .Y(n794) );
  INVX1 U69 ( .A(N14), .Y(n820) );
  INVX1 U71 ( .A(n501), .Y(n811) );
  INVX1 U72 ( .A(n502), .Y(n812) );
  INVX1 U73 ( .A(n503), .Y(n813) );
  INVX1 U75 ( .A(n504), .Y(n814) );
  INVX1 U77 ( .A(n505), .Y(n815) );
  INVX1 U79 ( .A(rst), .Y(n816) );
  INVX1 U81 ( .A(N12), .Y(n818) );
  INVX1 U83 ( .A(N13), .Y(n819) );
  INVX2 U84 ( .A(n794), .Y(n798) );
  INVX1 U85 ( .A(n801), .Y(n1) );
  INVX1 U87 ( .A(n1), .Y(n2) );
  INVX1 U89 ( .A(n817), .Y(n3) );
  INVX1 U91 ( .A(n801), .Y(n809) );
  MUX2X1 U93 ( .B(\mem<3><0> ), .A(\mem<2><0> ), .S(n799), .Y(n660) );
  INVX8 U95 ( .A(n790), .Y(n792) );
  INVX8 U96 ( .A(n793), .Y(n810) );
  MUX2X1 U97 ( .B(n651), .A(n650), .S(n793), .Y(n649) );
  MUX2X1 U99 ( .B(n657), .A(n656), .S(n793), .Y(n655) );
  MUX2X1 U101 ( .B(\mem<5><0> ), .A(\mem<4><0> ), .S(n2), .Y(n656) );
  MUX2X1 U103 ( .B(n660), .A(n659), .S(n793), .Y(n658) );
  MUX2X1 U105 ( .B(n747), .A(n746), .S(n793), .Y(n745) );
  MUX2X1 U107 ( .B(\mem<11><3> ), .A(\mem<10><3> ), .S(n799), .Y(n744) );
  MUX2X1 U108 ( .B(n752), .A(n753), .S(N13), .Y(n751) );
  MUX2X1 U109 ( .B(\mem<13><0> ), .A(\mem<12><0> ), .S(n801), .Y(n650) );
  MUX2X1 U111 ( .B(\mem<15><0> ), .A(\mem<14><0> ), .S(n799), .Y(n651) );
  MUX2X1 U113 ( .B(\mem<1><0> ), .A(\mem<0><0> ), .S(n801), .Y(n659) );
  MUX2X1 U115 ( .B(n649), .A(n652), .S(n790), .Y(n663) );
  AND2X2 U117 ( .A(N17), .B(n822), .Y(\data_out<4> ) );
  INVX1 U119 ( .A(n4), .Y(n5) );
  AND2X2 U120 ( .A(\mem<0><3> ), .B(n507), .Y(n6) );
  INVX1 U121 ( .A(n6), .Y(n7) );
  AND2X2 U123 ( .A(\mem<0><2> ), .B(n507), .Y(n8) );
  INVX1 U125 ( .A(n8), .Y(n9) );
  AND2X2 U127 ( .A(\mem<0><1> ), .B(n507), .Y(n10) );
  INVX1 U129 ( .A(n10), .Y(n11) );
  AND2X2 U131 ( .A(\mem<0><0> ), .B(n507), .Y(n12) );
  INVX1 U132 ( .A(n12), .Y(n13) );
  INVX1 U133 ( .A(n14), .Y(n15) );
  AND2X2 U135 ( .A(\mem<1><3> ), .B(n509), .Y(n16) );
  INVX1 U137 ( .A(n16), .Y(n17) );
  AND2X2 U139 ( .A(\mem<1><2> ), .B(n509), .Y(n18) );
  INVX1 U141 ( .A(n18), .Y(n19) );
  AND2X2 U143 ( .A(\mem<1><1> ), .B(n509), .Y(n20) );
  INVX1 U144 ( .A(n20), .Y(n21) );
  AND2X2 U145 ( .A(\mem<1><0> ), .B(n509), .Y(n22) );
  INVX1 U148 ( .A(n22), .Y(n23) );
  INVX1 U150 ( .A(n24), .Y(n25) );
  AND2X2 U152 ( .A(\mem<2><3> ), .B(n511), .Y(n26) );
  INVX1 U154 ( .A(n26), .Y(n27) );
  AND2X2 U156 ( .A(\mem<2><2> ), .B(n511), .Y(n28) );
  INVX1 U157 ( .A(n28), .Y(n29) );
  AND2X2 U158 ( .A(\mem<2><1> ), .B(n511), .Y(n30) );
  INVX1 U160 ( .A(n30), .Y(n31) );
  AND2X2 U162 ( .A(\mem<2><0> ), .B(n511), .Y(n32) );
  INVX1 U164 ( .A(n32), .Y(n33) );
  INVX1 U166 ( .A(n34), .Y(n35) );
  AND2X2 U168 ( .A(\mem<3><3> ), .B(n513), .Y(n36) );
  INVX1 U169 ( .A(n36), .Y(n37) );
  AND2X2 U170 ( .A(\mem<3><2> ), .B(n513), .Y(n38) );
  INVX1 U172 ( .A(n38), .Y(n39) );
  AND2X2 U174 ( .A(\mem<3><1> ), .B(n513), .Y(n40) );
  INVX1 U176 ( .A(n40), .Y(n41) );
  AND2X2 U178 ( .A(\mem<3><0> ), .B(n513), .Y(n42) );
  INVX1 U181 ( .A(n42), .Y(n43) );
  INVX1 U182 ( .A(n44), .Y(n45) );
  AND2X2 U184 ( .A(\mem<4><3> ), .B(n515), .Y(n46) );
  INVX1 U186 ( .A(n46), .Y(n47) );
  AND2X2 U188 ( .A(\mem<4><2> ), .B(n515), .Y(n48) );
  INVX1 U190 ( .A(n48), .Y(n49) );
  AND2X2 U192 ( .A(\mem<4><1> ), .B(n515), .Y(n50) );
  INVX1 U193 ( .A(n50), .Y(n51) );
  AND2X2 U194 ( .A(\mem<4><0> ), .B(n515), .Y(n52) );
  INVX1 U196 ( .A(n52), .Y(n53) );
  INVX1 U198 ( .A(n54), .Y(n55) );
  AND2X2 U200 ( .A(\mem<5><3> ), .B(n517), .Y(n58) );
  INVX1 U202 ( .A(n58), .Y(n59) );
  INVX1 U204 ( .A(n60), .Y(n61) );
  AND2X2 U205 ( .A(\mem<5><1> ), .B(n517), .Y(n62) );
  INVX1 U206 ( .A(n62), .Y(n63) );
  AND2X2 U208 ( .A(\mem<5><0> ), .B(n517), .Y(n64) );
  INVX1 U210 ( .A(n64), .Y(n66) );
  INVX1 U212 ( .A(n67), .Y(n68) );
  AND2X2 U214 ( .A(\mem<6><3> ), .B(n519), .Y(n69) );
  INVX1 U216 ( .A(n69), .Y(n70) );
  AND2X2 U217 ( .A(\mem<6><2> ), .B(n519), .Y(n71) );
  INVX1 U218 ( .A(n71), .Y(n72) );
  AND2X2 U220 ( .A(\mem<6><1> ), .B(n519), .Y(n74) );
  INVX1 U222 ( .A(n74), .Y(n75) );
  AND2X2 U224 ( .A(\mem<6><0> ), .B(n519), .Y(n76) );
  INVX1 U226 ( .A(n76), .Y(n77) );
  INVX1 U228 ( .A(n78), .Y(n79) );
  AND2X2 U229 ( .A(\mem<7><3> ), .B(n521), .Y(n80) );
  INVX1 U230 ( .A(n80), .Y(n82) );
  INVX1 U232 ( .A(n83), .Y(n84) );
  AND2X2 U234 ( .A(\mem<7><1> ), .B(n521), .Y(n85) );
  INVX1 U236 ( .A(n85), .Y(n86) );
  AND2X2 U238 ( .A(\mem<7><0> ), .B(n521), .Y(n87) );
  INVX1 U240 ( .A(n87), .Y(n88) );
  INVX1 U241 ( .A(n90), .Y(n91) );
  AND2X2 U242 ( .A(\mem<8><3> ), .B(n523), .Y(n92) );
  INVX1 U245 ( .A(n92), .Y(n93) );
  AND2X2 U247 ( .A(\mem<8><2> ), .B(n523), .Y(n94) );
  INVX1 U249 ( .A(n94), .Y(n95) );
  AND2X2 U251 ( .A(\mem<8><1> ), .B(n523), .Y(n96) );
  INVX1 U253 ( .A(n96), .Y(n98) );
  AND2X2 U254 ( .A(\mem<8><0> ), .B(n523), .Y(n99) );
  INVX1 U255 ( .A(n99), .Y(n100) );
  INVX1 U257 ( .A(n101), .Y(n102) );
  AND2X2 U259 ( .A(\mem<9><3> ), .B(n525), .Y(n103) );
  INVX1 U261 ( .A(n103), .Y(n104) );
  AND2X2 U263 ( .A(\mem<9><2> ), .B(n525), .Y(n106) );
  INVX1 U265 ( .A(n106), .Y(n107) );
  AND2X2 U266 ( .A(\mem<9><1> ), .B(n525), .Y(n108) );
  INVX1 U267 ( .A(n108), .Y(n109) );
  AND2X2 U269 ( .A(\mem<9><0> ), .B(n525), .Y(n110) );
  INVX1 U271 ( .A(n110), .Y(n111) );
  INVX1 U273 ( .A(n112), .Y(n116) );
  AND2X2 U275 ( .A(\mem<10><3> ), .B(n527), .Y(n117) );
  INVX1 U277 ( .A(n117), .Y(n118) );
  AND2X2 U278 ( .A(\mem<10><2> ), .B(n527), .Y(n119) );
  INVX1 U279 ( .A(n119), .Y(n120) );
  AND2X2 U281 ( .A(\mem<10><1> ), .B(n527), .Y(n121) );
  INVX1 U283 ( .A(n121), .Y(n122) );
  AND2X2 U285 ( .A(\mem<10><0> ), .B(n527), .Y(n123) );
  INVX1 U287 ( .A(n123), .Y(n124) );
  INVX1 U289 ( .A(n125), .Y(n126) );
  AND2X2 U290 ( .A(\mem<11><3> ), .B(n529), .Y(n127) );
  INVX1 U291 ( .A(n127), .Y(n128) );
  AND2X2 U293 ( .A(\mem<11><2> ), .B(n529), .Y(n129) );
  INVX1 U295 ( .A(n129), .Y(n130) );
  AND2X2 U297 ( .A(\mem<11><1> ), .B(n529), .Y(n131) );
  INVX1 U299 ( .A(n131), .Y(n132) );
  AND2X2 U301 ( .A(\mem<11><0> ), .B(n529), .Y(n133) );
  INVX1 U302 ( .A(n133), .Y(n134) );
  INVX1 U303 ( .A(n135), .Y(n137) );
  AND2X2 U305 ( .A(\mem<12><3> ), .B(n531), .Y(n138) );
  INVX1 U307 ( .A(n138), .Y(n139) );
  AND2X2 U309 ( .A(\mem<12><2> ), .B(n531), .Y(n140) );
  INVX1 U311 ( .A(n140), .Y(n141) );
  AND2X2 U313 ( .A(\mem<12><1> ), .B(n531), .Y(n142) );
  INVX1 U314 ( .A(n142), .Y(n143) );
  AND2X2 U315 ( .A(\mem<12><0> ), .B(n531), .Y(n144) );
  INVX1 U317 ( .A(n144), .Y(n145) );
  INVX1 U319 ( .A(n146), .Y(n147) );
  AND2X2 U321 ( .A(\mem<13><3> ), .B(n533), .Y(n148) );
  INVX1 U323 ( .A(n148), .Y(n149) );
  INVX1 U325 ( .A(n150), .Y(n151) );
  AND2X2 U326 ( .A(\mem<13><1> ), .B(n533), .Y(n152) );
  INVX1 U327 ( .A(n152), .Y(n153) );
  AND2X2 U329 ( .A(\mem<13><0> ), .B(n533), .Y(n154) );
  INVX1 U331 ( .A(n154), .Y(n155) );
  INVX1 U333 ( .A(n156), .Y(n157) );
  AND2X2 U335 ( .A(\mem<14><3> ), .B(n535), .Y(n158) );
  INVX1 U337 ( .A(n158), .Y(n159) );
  AND2X2 U338 ( .A(\mem<14><2> ), .B(n535), .Y(n160) );
  INVX1 U339 ( .A(n160), .Y(n161) );
  AND2X2 U342 ( .A(\mem<14><1> ), .B(n535), .Y(n162) );
  INVX1 U344 ( .A(n162), .Y(n163) );
  AND2X2 U346 ( .A(\mem<14><0> ), .B(n535), .Y(n164) );
  INVX1 U348 ( .A(n164), .Y(n165) );
  INVX1 U350 ( .A(n166), .Y(n167) );
  AND2X2 U351 ( .A(\mem<15><3> ), .B(n537), .Y(n168) );
  INVX1 U352 ( .A(n168), .Y(n169) );
  INVX1 U355 ( .A(n170), .Y(n171) );
  AND2X2 U357 ( .A(\mem<15><1> ), .B(n537), .Y(n173) );
  INVX1 U359 ( .A(n173), .Y(n174) );
  AND2X2 U361 ( .A(\mem<15><0> ), .B(n537), .Y(n175) );
  INVX1 U363 ( .A(n175), .Y(n176) );
  INVX1 U364 ( .A(n177), .Y(n178) );
  AND2X2 U365 ( .A(\mem<16><3> ), .B(n539), .Y(n179) );
  INVX1 U368 ( .A(n179), .Y(n180) );
  AND2X2 U370 ( .A(\mem<16><2> ), .B(n539), .Y(n181) );
  INVX1 U372 ( .A(n181), .Y(n182) );
  AND2X2 U374 ( .A(\mem<16><1> ), .B(n539), .Y(n183) );
  INVX1 U376 ( .A(n183), .Y(n184) );
  AND2X2 U377 ( .A(\mem<16><0> ), .B(n539), .Y(n185) );
  INVX1 U378 ( .A(n185), .Y(n186) );
  INVX1 U381 ( .A(n187), .Y(n188) );
  AND2X2 U383 ( .A(\mem<17><3> ), .B(n541), .Y(n189) );
  INVX1 U385 ( .A(n189), .Y(n190) );
  INVX1 U387 ( .A(n191), .Y(n192) );
  AND2X2 U389 ( .A(\mem<17><1> ), .B(n541), .Y(n193) );
  INVX1 U390 ( .A(n193), .Y(n194) );
  AND2X2 U391 ( .A(\mem<17><0> ), .B(n541), .Y(n195) );
  INVX1 U394 ( .A(n195), .Y(n196) );
  INVX1 U396 ( .A(n197), .Y(n198) );
  AND2X2 U398 ( .A(\mem<18><3> ), .B(n543), .Y(n199) );
  INVX1 U400 ( .A(n199), .Y(n200) );
  AND2X2 U402 ( .A(\mem<18><2> ), .B(n543), .Y(n201) );
  INVX1 U403 ( .A(n201), .Y(n202) );
  AND2X2 U404 ( .A(\mem<18><1> ), .B(n543), .Y(n203) );
  INVX1 U407 ( .A(n203), .Y(n204) );
  AND2X2 U409 ( .A(\mem<18><0> ), .B(n543), .Y(n205) );
  INVX1 U411 ( .A(n205), .Y(n206) );
  INVX1 U413 ( .A(n207), .Y(n208) );
  AND2X2 U415 ( .A(\mem<19><3> ), .B(n545), .Y(n209) );
  INVX1 U416 ( .A(n209), .Y(n210) );
  INVX1 U417 ( .A(n211), .Y(n212) );
  AND2X2 U420 ( .A(\mem<19><1> ), .B(n545), .Y(n213) );
  INVX1 U422 ( .A(n213), .Y(n214) );
  AND2X2 U424 ( .A(\mem<19><0> ), .B(n545), .Y(n215) );
  INVX1 U426 ( .A(n215), .Y(n216) );
  INVX1 U428 ( .A(n217), .Y(n218) );
  AND2X2 U429 ( .A(\mem<20><3> ), .B(n547), .Y(n219) );
  INVX1 U430 ( .A(n219), .Y(n220) );
  INVX1 U433 ( .A(n221), .Y(n222) );
  AND2X2 U434 ( .A(\mem<20><1> ), .B(n547), .Y(n223) );
  INVX1 U436 ( .A(n223), .Y(n224) );
  AND2X2 U437 ( .A(\mem<20><0> ), .B(n547), .Y(n225) );
  INVX1 U439 ( .A(n225), .Y(n226) );
  INVX1 U440 ( .A(n227), .Y(n228) );
  INVX1 U442 ( .A(n230), .Y(n231) );
  INVX1 U443 ( .A(n232), .Y(n233) );
  AND2X2 U445 ( .A(\mem<21><0> ), .B(n549), .Y(n234) );
  INVX1 U446 ( .A(n234), .Y(n235) );
  INVX1 U447 ( .A(n236), .Y(n237) );
  AND2X2 U451 ( .A(\mem<22><3> ), .B(n551), .Y(n238) );
  INVX1 U452 ( .A(n238), .Y(n239) );
  INVX1 U453 ( .A(n240), .Y(n241) );
  AND2X2 U454 ( .A(\mem<22><1> ), .B(n551), .Y(n242) );
  INVX1 U455 ( .A(n242), .Y(n243) );
  AND2X2 U456 ( .A(\mem<22><0> ), .B(n551), .Y(n244) );
  INVX1 U457 ( .A(n244), .Y(n245) );
  INVX1 U458 ( .A(n246), .Y(n247) );
  INVX1 U459 ( .A(n248), .Y(n249) );
  INVX1 U460 ( .A(n250), .Y(n251) );
  INVX1 U461 ( .A(n252), .Y(n253) );
  AND2X2 U462 ( .A(\mem<23><0> ), .B(n553), .Y(n254) );
  INVX1 U463 ( .A(n254), .Y(n255) );
  INVX1 U464 ( .A(n256), .Y(n257) );
  AND2X2 U465 ( .A(\mem<24><3> ), .B(n555), .Y(n258) );
  INVX1 U466 ( .A(n258), .Y(n259) );
  AND2X2 U467 ( .A(\mem<24><2> ), .B(n555), .Y(n260) );
  INVX1 U468 ( .A(n260), .Y(n261) );
  AND2X2 U469 ( .A(\mem<24><1> ), .B(n555), .Y(n262) );
  INVX1 U470 ( .A(n262), .Y(n263) );
  AND2X2 U471 ( .A(\mem<24><0> ), .B(n555), .Y(n264) );
  INVX1 U472 ( .A(n264), .Y(n265) );
  INVX1 U473 ( .A(n266), .Y(n267) );
  AND2X2 U474 ( .A(\mem<25><3> ), .B(n557), .Y(n268) );
  INVX1 U475 ( .A(n268), .Y(n269) );
  INVX1 U476 ( .A(n270), .Y(n271) );
  AND2X2 U477 ( .A(\mem<25><1> ), .B(n557), .Y(n272) );
  INVX1 U478 ( .A(n272), .Y(n273) );
  AND2X2 U479 ( .A(\mem<25><0> ), .B(n557), .Y(n274) );
  INVX1 U480 ( .A(n274), .Y(n275) );
  INVX1 U481 ( .A(n276), .Y(n277) );
  AND2X2 U482 ( .A(\mem<26><3> ), .B(n559), .Y(n278) );
  INVX1 U483 ( .A(n278), .Y(n279) );
  AND2X2 U484 ( .A(\mem<26><2> ), .B(n559), .Y(n280) );
  INVX1 U485 ( .A(n280), .Y(n281) );
  AND2X2 U486 ( .A(\mem<26><1> ), .B(n559), .Y(n282) );
  INVX1 U487 ( .A(n282), .Y(n283) );
  AND2X2 U488 ( .A(\mem<26><0> ), .B(n559), .Y(n284) );
  INVX1 U489 ( .A(n284), .Y(n285) );
  INVX1 U490 ( .A(n287), .Y(n448) );
  AND2X2 U491 ( .A(\mem<27><3> ), .B(n561), .Y(n449) );
  INVX1 U492 ( .A(n449), .Y(n450) );
  INVX1 U493 ( .A(n451), .Y(n452) );
  AND2X2 U494 ( .A(\mem<27><1> ), .B(n561), .Y(n453) );
  INVX1 U495 ( .A(n453), .Y(n454) );
  AND2X2 U496 ( .A(\mem<27><0> ), .B(n561), .Y(n455) );
  INVX1 U497 ( .A(n455), .Y(n456) );
  INVX1 U498 ( .A(n457), .Y(n458) );
  AND2X2 U499 ( .A(\mem<28><3> ), .B(n563), .Y(n459) );
  INVX1 U500 ( .A(n459), .Y(n460) );
  INVX1 U501 ( .A(n461), .Y(n462) );
  AND2X2 U502 ( .A(\mem<28><1> ), .B(n563), .Y(n463) );
  INVX1 U503 ( .A(n463), .Y(n464) );
  AND2X2 U504 ( .A(\mem<28><0> ), .B(n563), .Y(n465) );
  INVX1 U505 ( .A(n465), .Y(n466) );
  INVX1 U506 ( .A(n467), .Y(n468) );
  INVX1 U507 ( .A(n469), .Y(n470) );
  INVX1 U508 ( .A(n471), .Y(n472) );
  INVX1 U509 ( .A(n473), .Y(n474) );
  AND2X2 U510 ( .A(\mem<29><0> ), .B(n565), .Y(n475) );
  INVX1 U511 ( .A(n475), .Y(n476) );
  INVX1 U512 ( .A(n477), .Y(n478) );
  AND2X2 U513 ( .A(\mem<30><3> ), .B(n567), .Y(n479) );
  INVX1 U514 ( .A(n479), .Y(n480) );
  INVX1 U515 ( .A(n481), .Y(n482) );
  AND2X2 U516 ( .A(\mem<30><1> ), .B(n567), .Y(n483) );
  INVX1 U517 ( .A(n483), .Y(n484) );
  AND2X2 U518 ( .A(\mem<30><0> ), .B(n567), .Y(n485) );
  INVX1 U519 ( .A(n485), .Y(n486) );
  INVX1 U520 ( .A(n487), .Y(n488) );
  INVX1 U521 ( .A(n489), .Y(n490) );
  INVX1 U522 ( .A(n491), .Y(n492) );
  INVX1 U523 ( .A(n493), .Y(n494) );
  AND2X2 U524 ( .A(\mem<31><0> ), .B(n569), .Y(n495) );
  INVX1 U525 ( .A(n495), .Y(n496) );
  BUFX2 U526 ( .A(n286), .Y(n497) );
  INVX1 U527 ( .A(n497), .Y(n823) );
  BUFX2 U528 ( .A(n229), .Y(n498) );
  INVX1 U529 ( .A(n498), .Y(n824) );
  BUFX2 U530 ( .A(n172), .Y(n499) );
  INVX1 U531 ( .A(n499), .Y(n825) );
  BUFX2 U532 ( .A(n114), .Y(n500) );
  INVX1 U533 ( .A(n500), .Y(n826) );
  AND2X1 U534 ( .A(\data_in<4> ), .B(n56), .Y(n501) );
  AND2X1 U535 ( .A(\data_in<3> ), .B(n56), .Y(n502) );
  AND2X1 U536 ( .A(\data_in<2> ), .B(n56), .Y(n503) );
  AND2X1 U537 ( .A(\data_in<1> ), .B(n56), .Y(n504) );
  AND2X1 U538 ( .A(\data_in<0> ), .B(n56), .Y(n505) );
  AND2X1 U539 ( .A(n572), .B(n56), .Y(n506) );
  INVX1 U540 ( .A(n506), .Y(n507) );
  AND2X1 U541 ( .A(n574), .B(n56), .Y(n508) );
  INVX1 U542 ( .A(n508), .Y(n509) );
  AND2X1 U543 ( .A(n576), .B(n56), .Y(n510) );
  INVX1 U544 ( .A(n510), .Y(n511) );
  AND2X1 U545 ( .A(n578), .B(n56), .Y(n512) );
  INVX1 U546 ( .A(n512), .Y(n513) );
  AND2X1 U547 ( .A(n580), .B(n56), .Y(n514) );
  INVX1 U548 ( .A(n514), .Y(n515) );
  AND2X1 U549 ( .A(n582), .B(n56), .Y(n516) );
  INVX1 U550 ( .A(n516), .Y(n517) );
  AND2X1 U551 ( .A(n584), .B(n56), .Y(n518) );
  INVX1 U552 ( .A(n518), .Y(n519) );
  AND2X1 U553 ( .A(n586), .B(n56), .Y(n520) );
  INVX1 U554 ( .A(n520), .Y(n521) );
  AND2X1 U555 ( .A(n588), .B(n56), .Y(n522) );
  INVX1 U556 ( .A(n522), .Y(n523) );
  AND2X1 U557 ( .A(n590), .B(n56), .Y(n524) );
  INVX1 U558 ( .A(n524), .Y(n525) );
  AND2X1 U559 ( .A(n592), .B(n56), .Y(n526) );
  INVX1 U560 ( .A(n526), .Y(n527) );
  AND2X1 U561 ( .A(n594), .B(n56), .Y(n528) );
  INVX1 U562 ( .A(n528), .Y(n529) );
  AND2X1 U563 ( .A(n596), .B(n56), .Y(n530) );
  INVX1 U564 ( .A(n530), .Y(n531) );
  AND2X1 U565 ( .A(n598), .B(n56), .Y(n532) );
  INVX1 U566 ( .A(n532), .Y(n533) );
  AND2X1 U567 ( .A(n600), .B(n56), .Y(n534) );
  INVX1 U568 ( .A(n534), .Y(n535) );
  AND2X1 U569 ( .A(n602), .B(n56), .Y(n536) );
  INVX1 U570 ( .A(n536), .Y(n537) );
  AND2X1 U571 ( .A(n604), .B(n56), .Y(n538) );
  INVX1 U572 ( .A(n538), .Y(n539) );
  AND2X1 U573 ( .A(n606), .B(n56), .Y(n540) );
  INVX1 U574 ( .A(n540), .Y(n541) );
  AND2X1 U575 ( .A(n608), .B(n56), .Y(n542) );
  INVX1 U576 ( .A(n542), .Y(n543) );
  AND2X1 U577 ( .A(n610), .B(n56), .Y(n544) );
  INVX1 U578 ( .A(n544), .Y(n545) );
  AND2X1 U579 ( .A(n612), .B(n56), .Y(n546) );
  INVX1 U580 ( .A(n546), .Y(n547) );
  AND2X1 U581 ( .A(n614), .B(n56), .Y(n548) );
  INVX1 U582 ( .A(n548), .Y(n549) );
  AND2X1 U583 ( .A(n616), .B(n56), .Y(n550) );
  INVX1 U584 ( .A(n550), .Y(n551) );
  AND2X1 U585 ( .A(n618), .B(n56), .Y(n552) );
  INVX1 U586 ( .A(n552), .Y(n553) );
  AND2X1 U587 ( .A(n620), .B(n56), .Y(n554) );
  INVX1 U588 ( .A(n554), .Y(n555) );
  AND2X1 U589 ( .A(n622), .B(n56), .Y(n556) );
  INVX1 U590 ( .A(n556), .Y(n557) );
  AND2X1 U591 ( .A(n624), .B(n56), .Y(n558) );
  INVX1 U592 ( .A(n558), .Y(n559) );
  AND2X1 U593 ( .A(n626), .B(n56), .Y(n560) );
  INVX1 U594 ( .A(n560), .Y(n561) );
  AND2X1 U595 ( .A(n628), .B(n56), .Y(n562) );
  INVX1 U596 ( .A(n562), .Y(n563) );
  AND2X1 U597 ( .A(n630), .B(n56), .Y(n564) );
  INVX1 U598 ( .A(n564), .Y(n565) );
  AND2X1 U599 ( .A(n632), .B(n56), .Y(n566) );
  INVX1 U600 ( .A(n566), .Y(n567) );
  AND2X1 U601 ( .A(n570), .B(n56), .Y(n568) );
  INVX1 U602 ( .A(n568), .Y(n569) );
  AND2X1 U603 ( .A(n57), .B(n826), .Y(n570) );
  INVX1 U604 ( .A(n570), .Y(n571) );
  AND2X1 U605 ( .A(n823), .B(n113), .Y(n572) );
  INVX1 U606 ( .A(n572), .Y(n573) );
  AND2X1 U607 ( .A(n823), .B(n105), .Y(n574) );
  INVX1 U608 ( .A(n574), .Y(n575) );
  AND2X1 U609 ( .A(n823), .B(n97), .Y(n576) );
  INVX1 U610 ( .A(n576), .Y(n577) );
  AND2X1 U611 ( .A(n823), .B(n89), .Y(n578) );
  INVX1 U612 ( .A(n578), .Y(n579) );
  AND2X1 U613 ( .A(n823), .B(n81), .Y(n580) );
  INVX1 U614 ( .A(n580), .Y(n581) );
  AND2X1 U615 ( .A(n823), .B(n73), .Y(n582) );
  INVX1 U616 ( .A(n582), .Y(n583) );
  AND2X1 U617 ( .A(n823), .B(n65), .Y(n584) );
  INVX1 U618 ( .A(n584), .Y(n585) );
  AND2X1 U619 ( .A(n823), .B(n57), .Y(n586) );
  INVX1 U620 ( .A(n586), .Y(n587) );
  AND2X1 U621 ( .A(n824), .B(n113), .Y(n588) );
  INVX1 U622 ( .A(n588), .Y(n589) );
  AND2X1 U623 ( .A(n824), .B(n105), .Y(n590) );
  INVX1 U624 ( .A(n590), .Y(n591) );
  AND2X1 U625 ( .A(n824), .B(n97), .Y(n592) );
  INVX1 U626 ( .A(n592), .Y(n593) );
  AND2X1 U627 ( .A(n824), .B(n89), .Y(n594) );
  INVX1 U628 ( .A(n594), .Y(n595) );
  AND2X1 U629 ( .A(n824), .B(n81), .Y(n596) );
  INVX1 U630 ( .A(n596), .Y(n597) );
  AND2X1 U631 ( .A(n824), .B(n73), .Y(n598) );
  INVX1 U632 ( .A(n598), .Y(n599) );
  AND2X1 U633 ( .A(n824), .B(n65), .Y(n600) );
  INVX1 U634 ( .A(n600), .Y(n601) );
  AND2X1 U635 ( .A(n824), .B(n57), .Y(n602) );
  INVX1 U636 ( .A(n602), .Y(n603) );
  AND2X1 U637 ( .A(n825), .B(n113), .Y(n604) );
  INVX1 U638 ( .A(n604), .Y(n605) );
  AND2X1 U639 ( .A(n825), .B(n105), .Y(n606) );
  INVX1 U640 ( .A(n606), .Y(n607) );
  AND2X1 U641 ( .A(n825), .B(n97), .Y(n608) );
  INVX1 U642 ( .A(n608), .Y(n609) );
  AND2X1 U643 ( .A(n825), .B(n89), .Y(n610) );
  INVX1 U644 ( .A(n610), .Y(n611) );
  AND2X1 U645 ( .A(n825), .B(n81), .Y(n612) );
  INVX1 U646 ( .A(n612), .Y(n613) );
  AND2X1 U647 ( .A(n825), .B(n73), .Y(n614) );
  INVX1 U648 ( .A(n614), .Y(n615) );
  AND2X1 U649 ( .A(n825), .B(n65), .Y(n616) );
  INVX1 U650 ( .A(n616), .Y(n617) );
  AND2X1 U651 ( .A(n825), .B(n57), .Y(n618) );
  INVX1 U652 ( .A(n618), .Y(n619) );
  AND2X1 U653 ( .A(n113), .B(n826), .Y(n620) );
  INVX1 U654 ( .A(n620), .Y(n621) );
  AND2X1 U655 ( .A(n105), .B(n826), .Y(n622) );
  INVX1 U656 ( .A(n622), .Y(n623) );
  AND2X1 U657 ( .A(n97), .B(n826), .Y(n624) );
  INVX1 U658 ( .A(n624), .Y(n625) );
  AND2X1 U659 ( .A(n89), .B(n826), .Y(n626) );
  INVX1 U660 ( .A(n626), .Y(n627) );
  AND2X1 U661 ( .A(n81), .B(n826), .Y(n628) );
  INVX1 U662 ( .A(n628), .Y(n629) );
  AND2X1 U663 ( .A(n73), .B(n826), .Y(n630) );
  INVX1 U664 ( .A(n630), .Y(n631) );
  AND2X1 U665 ( .A(n65), .B(n826), .Y(n632) );
  INVX1 U666 ( .A(n632), .Y(n633) );
  MUX2X1 U667 ( .B(n635), .A(n636), .S(n810), .Y(n634) );
  MUX2X1 U668 ( .B(n638), .A(n639), .S(n798), .Y(n637) );
  MUX2X1 U669 ( .B(n641), .A(n642), .S(n810), .Y(n640) );
  MUX2X1 U670 ( .B(n644), .A(n645), .S(n798), .Y(n643) );
  MUX2X1 U671 ( .B(n647), .A(n648), .S(n789), .Y(n646) );
  MUX2X1 U672 ( .B(n653), .A(n654), .S(n798), .Y(n652) );
  MUX2X1 U673 ( .B(n662), .A(n663), .S(n789), .Y(n661) );
  MUX2X1 U674 ( .B(n665), .A(n666), .S(n810), .Y(n664) );
  MUX2X1 U675 ( .B(n668), .A(n669), .S(n798), .Y(n667) );
  MUX2X1 U676 ( .B(n671), .A(n672), .S(n810), .Y(n670) );
  MUX2X1 U677 ( .B(n674), .A(n675), .S(n798), .Y(n673) );
  MUX2X1 U678 ( .B(n677), .A(n678), .S(n789), .Y(n676) );
  MUX2X1 U679 ( .B(n680), .A(n681), .S(n795), .Y(n679) );
  MUX2X1 U680 ( .B(n683), .A(n684), .S(n797), .Y(n682) );
  MUX2X1 U681 ( .B(n686), .A(n687), .S(n795), .Y(n685) );
  MUX2X1 U682 ( .B(n689), .A(n690), .S(n797), .Y(n688) );
  MUX2X1 U683 ( .B(n692), .A(n693), .S(n789), .Y(n691) );
  MUX2X1 U684 ( .B(n695), .A(n696), .S(n796), .Y(n694) );
  MUX2X1 U685 ( .B(n698), .A(n699), .S(n796), .Y(n697) );
  MUX2X1 U686 ( .B(n701), .A(n702), .S(n796), .Y(n700) );
  MUX2X1 U687 ( .B(n704), .A(n705), .S(n796), .Y(n703) );
  MUX2X1 U688 ( .B(n707), .A(n708), .S(n789), .Y(n706) );
  MUX2X1 U689 ( .B(n710), .A(n711), .S(n795), .Y(n709) );
  MUX2X1 U690 ( .B(n713), .A(n714), .S(n797), .Y(n712) );
  MUX2X1 U691 ( .B(n716), .A(n717), .S(n796), .Y(n715) );
  MUX2X1 U692 ( .B(n719), .A(n720), .S(n797), .Y(n718) );
  MUX2X1 U693 ( .B(n722), .A(n723), .S(n789), .Y(n721) );
  MUX2X1 U694 ( .B(n725), .A(n726), .S(n795), .Y(n724) );
  MUX2X1 U695 ( .B(n728), .A(n729), .S(n795), .Y(n727) );
  MUX2X1 U696 ( .B(n731), .A(n732), .S(n796), .Y(n730) );
  MUX2X1 U697 ( .B(n734), .A(n735), .S(n795), .Y(n733) );
  MUX2X1 U698 ( .B(n737), .A(n738), .S(n789), .Y(n736) );
  MUX2X1 U699 ( .B(n740), .A(n741), .S(n795), .Y(n739) );
  MUX2X1 U700 ( .B(n743), .A(n744), .S(n797), .Y(n742) );
  MUX2X1 U701 ( .B(n749), .A(n750), .S(n797), .Y(n748) );
  MUX2X1 U702 ( .B(n755), .A(n756), .S(n796), .Y(n754) );
  MUX2X1 U703 ( .B(n758), .A(n759), .S(n796), .Y(n757) );
  MUX2X1 U704 ( .B(n761), .A(n762), .S(n797), .Y(n760) );
  MUX2X1 U705 ( .B(n764), .A(n765), .S(n796), .Y(n763) );
  MUX2X1 U706 ( .B(n767), .A(n768), .S(n789), .Y(n766) );
  MUX2X1 U707 ( .B(n770), .A(n771), .S(n796), .Y(n769) );
  MUX2X1 U708 ( .B(n773), .A(n774), .S(n796), .Y(n772) );
  MUX2X1 U709 ( .B(n776), .A(n777), .S(n796), .Y(n775) );
  MUX2X1 U710 ( .B(n779), .A(n780), .S(n796), .Y(n778) );
  MUX2X1 U711 ( .B(n782), .A(n783), .S(n789), .Y(n781) );
  MUX2X1 U712 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n805), .Y(n636) );
  MUX2X1 U713 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n807), .Y(n635) );
  MUX2X1 U714 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n808), .Y(n639) );
  MUX2X1 U715 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n808), .Y(n638) );
  MUX2X1 U716 ( .B(n637), .A(n634), .S(n792), .Y(n648) );
  MUX2X1 U717 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n804), .Y(n642) );
  MUX2X1 U718 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n802), .Y(n641) );
  MUX2X1 U719 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n808), .Y(n645) );
  MUX2X1 U720 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n805), .Y(n644) );
  MUX2X1 U721 ( .B(n643), .A(n640), .S(n791), .Y(n647) );
  MUX2X1 U722 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n808), .Y(n654) );
  MUX2X1 U723 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n808), .Y(n653) );
  MUX2X1 U724 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n807), .Y(n657) );
  MUX2X1 U725 ( .B(n658), .A(n655), .S(n792), .Y(n662) );
  MUX2X1 U726 ( .B(n661), .A(n646), .S(N14), .Y(n784) );
  MUX2X1 U727 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n806), .Y(n666) );
  MUX2X1 U728 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n807), .Y(n665) );
  MUX2X1 U729 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n806), .Y(n669) );
  MUX2X1 U730 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n806), .Y(n668) );
  MUX2X1 U731 ( .B(n667), .A(n664), .S(n791), .Y(n678) );
  MUX2X1 U732 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n802), .Y(n672) );
  MUX2X1 U733 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n806), .Y(n671) );
  MUX2X1 U734 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n807), .Y(n675) );
  MUX2X1 U735 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n806), .Y(n674) );
  MUX2X1 U736 ( .B(n673), .A(n670), .S(n791), .Y(n677) );
  MUX2X1 U737 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n807), .Y(n681) );
  MUX2X1 U738 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n806), .Y(n680) );
  MUX2X1 U739 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n808), .Y(n684) );
  MUX2X1 U740 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n805), .Y(n683) );
  MUX2X1 U741 ( .B(n682), .A(n679), .S(n792), .Y(n693) );
  MUX2X1 U742 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n805), .Y(n687) );
  MUX2X1 U743 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n805), .Y(n686) );
  MUX2X1 U744 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n807), .Y(n690) );
  MUX2X1 U745 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n807), .Y(n689) );
  MUX2X1 U746 ( .B(n688), .A(n685), .S(n792), .Y(n692) );
  MUX2X1 U747 ( .B(n691), .A(n676), .S(N14), .Y(n785) );
  MUX2X1 U748 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n807), .Y(n696) );
  MUX2X1 U749 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n805), .Y(n695) );
  MUX2X1 U750 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n805), .Y(n699) );
  MUX2X1 U751 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n806), .Y(n698) );
  MUX2X1 U752 ( .B(n697), .A(n694), .S(n791), .Y(n708) );
  MUX2X1 U753 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n806), .Y(n702) );
  MUX2X1 U754 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n802), .Y(n701) );
  MUX2X1 U755 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n806), .Y(n705) );
  MUX2X1 U756 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n806), .Y(n704) );
  MUX2X1 U757 ( .B(n703), .A(n700), .S(n791), .Y(n707) );
  MUX2X1 U758 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n806), .Y(n711) );
  MUX2X1 U759 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n807), .Y(n710) );
  MUX2X1 U760 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n805), .Y(n714) );
  MUX2X1 U761 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n807), .Y(n713) );
  MUX2X1 U762 ( .B(n712), .A(n709), .S(n791), .Y(n723) );
  MUX2X1 U763 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n805), .Y(n717) );
  MUX2X1 U764 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n805), .Y(n716) );
  MUX2X1 U765 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n805), .Y(n720) );
  MUX2X1 U766 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n807), .Y(n719) );
  MUX2X1 U767 ( .B(n718), .A(n715), .S(n791), .Y(n722) );
  MUX2X1 U768 ( .B(n721), .A(n706), .S(N14), .Y(n786) );
  MUX2X1 U769 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n803), .Y(n726) );
  MUX2X1 U770 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n803), .Y(n725) );
  MUX2X1 U771 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n804), .Y(n729) );
  MUX2X1 U772 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n804), .Y(n728) );
  MUX2X1 U773 ( .B(n727), .A(n724), .S(n791), .Y(n738) );
  MUX2X1 U774 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n802), .Y(n732) );
  MUX2X1 U775 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n809), .Y(n731) );
  MUX2X1 U776 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n803), .Y(n735) );
  MUX2X1 U777 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n803), .Y(n734) );
  MUX2X1 U778 ( .B(n733), .A(n730), .S(n791), .Y(n737) );
  MUX2X1 U779 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n804), .Y(n741) );
  MUX2X1 U780 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n803), .Y(n740) );
  MUX2X1 U781 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n804), .Y(n743) );
  MUX2X1 U782 ( .B(n742), .A(n739), .S(n792), .Y(n753) );
  MUX2X1 U783 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n802), .Y(n747) );
  MUX2X1 U784 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n802), .Y(n746) );
  MUX2X1 U785 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n808), .Y(n750) );
  MUX2X1 U786 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n804), .Y(n749) );
  MUX2X1 U787 ( .B(n748), .A(n745), .S(n792), .Y(n752) );
  MUX2X1 U788 ( .B(n751), .A(n736), .S(N14), .Y(n787) );
  MUX2X1 U789 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n802), .Y(n756) );
  MUX2X1 U790 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n803), .Y(n755) );
  MUX2X1 U791 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n803), .Y(n759) );
  MUX2X1 U792 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n809), .Y(n758) );
  MUX2X1 U793 ( .B(n757), .A(n754), .S(n791), .Y(n768) );
  MUX2X1 U794 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n802), .Y(n762) );
  MUX2X1 U795 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n803), .Y(n761) );
  MUX2X1 U796 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n802), .Y(n765) );
  MUX2X1 U797 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n803), .Y(n764) );
  MUX2X1 U798 ( .B(n763), .A(n760), .S(n791), .Y(n767) );
  MUX2X1 U799 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n802), .Y(n771) );
  MUX2X1 U800 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n802), .Y(n770) );
  MUX2X1 U801 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n803), .Y(n774) );
  MUX2X1 U802 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n802), .Y(n773) );
  MUX2X1 U803 ( .B(n772), .A(n769), .S(n791), .Y(n783) );
  MUX2X1 U804 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n803), .Y(n777) );
  MUX2X1 U805 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n802), .Y(n776) );
  MUX2X1 U806 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n803), .Y(n780) );
  MUX2X1 U807 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n803), .Y(n779) );
  MUX2X1 U808 ( .B(n778), .A(n775), .S(n791), .Y(n782) );
  MUX2X1 U809 ( .B(n781), .A(n766), .S(N14), .Y(n788) );
  INVX8 U810 ( .A(n819), .Y(n789) );
  INVX8 U811 ( .A(N12), .Y(n790) );
  INVX8 U812 ( .A(n790), .Y(n791) );
  INVX8 U813 ( .A(n794), .Y(n795) );
  INVX8 U814 ( .A(n794), .Y(n796) );
  INVX8 U815 ( .A(n793), .Y(n797) );
  INVX8 U816 ( .A(N10), .Y(n800) );
  INVX8 U817 ( .A(N10), .Y(n801) );
  INVX8 U818 ( .A(n801), .Y(n802) );
  INVX8 U819 ( .A(n801), .Y(n803) );
  INVX8 U820 ( .A(n801), .Y(n804) );
  INVX8 U821 ( .A(n800), .Y(n805) );
  INVX8 U822 ( .A(n799), .Y(n806) );
  INVX8 U823 ( .A(n800), .Y(n807) );
  INVX8 U824 ( .A(n800), .Y(n808) );
  INVX1 U825 ( .A(n786), .Y(N19) );
  INVX1 U826 ( .A(n787), .Y(N18) );
  INVX1 U827 ( .A(n785), .Y(N20) );
  INVX1 U828 ( .A(n784), .Y(N21) );
  INVX4 U829 ( .A(N10), .Y(n799) );
  INVX4 U830 ( .A(N11), .Y(n793) );
  INVX1 U831 ( .A(n809), .Y(n817) );
  OR2X2 U832 ( .A(write), .B(rst), .Y(n821) );
  INVX2 U833 ( .A(n821), .Y(n822) );
  AND2X2 U834 ( .A(N21), .B(n822), .Y(\data_out<0> ) );
  AND2X2 U835 ( .A(N20), .B(n822), .Y(\data_out<1> ) );
  AND2X2 U836 ( .A(N19), .B(n822), .Y(\data_out<2> ) );
  AND2X2 U837 ( .A(N18), .B(n822), .Y(\data_out<3> ) );
endmodule


module memc_Size1 ( .data_out(\data_out<0> ), .addr({\addr<7> , \addr<6> , 
        \addr<5> , \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), 
    .data_in(\data_in<0> ), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<0> , write, clk, rst, createdump,
         \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> ;
  output \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><0> , \mem<1><0> , \mem<2><0> ,
         \mem<3><0> , \mem<4><0> , \mem<5><0> , \mem<6><0> , \mem<7><0> ,
         \mem<8><0> , \mem<9><0> , \mem<10><0> , \mem<11><0> , \mem<12><0> ,
         \mem<13><0> , \mem<14><0> , \mem<15><0> , \mem<16><0> , \mem<17><0> ,
         \mem<18><0> , \mem<19><0> , \mem<20><0> , \mem<21><0> , \mem<22><0> ,
         \mem<23><0> , \mem<24><0> , \mem<25><0> , \mem<26><0> , \mem<27><0> ,
         \mem<28><0> , \mem<29><0> , \mem<30><0> , \mem<31><0> , n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><0>  ( .D(n92), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n91), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n90), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n89), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n88), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n87), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n86), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n85), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n84), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n83), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n82), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n81), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n80), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n79), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n78), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n77), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n76), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n75), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n74), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n73), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n72), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n71), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n70), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n69), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n68), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n67), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n66), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n65), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n64), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n63), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n62), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n61), .CLK(clk), .Q(\mem<31><0> ) );
  NOR3X1 U93 ( .A(n158), .B(n2), .C(n150), .Y(\data_out<0> ) );
  INVX1 U2 ( .A(n163), .Y(n151) );
  INVX1 U3 ( .A(n159), .Y(n158) );
  AND2X1 U4 ( .A(n116), .B(n57), .Y(n36) );
  AND2X1 U5 ( .A(n113), .B(n57), .Y(n38) );
  AND2X1 U6 ( .A(n97), .B(n57), .Y(n40) );
  AND2X1 U7 ( .A(n100), .B(n57), .Y(n42) );
  AND2X1 U8 ( .A(n103), .B(n57), .Y(n44) );
  AND2X1 U9 ( .A(n106), .B(n57), .Y(n46) );
  AND2X1 U10 ( .A(n109), .B(n57), .Y(n48) );
  AND2X1 U11 ( .A(n115), .B(n57), .Y(n50) );
  AND2X1 U12 ( .A(n161), .B(n93), .Y(n115) );
  INVX2 U13 ( .A(n155), .Y(n156) );
  INVX2 U14 ( .A(n153), .Y(n154) );
  INVX1 U15 ( .A(n161), .Y(n152) );
  NOR3X1 U16 ( .A(n95), .B(n167), .C(N14), .Y(n1) );
  INVX2 U17 ( .A(n1), .Y(n195) );
  INVX1 U18 ( .A(N14), .Y(n169) );
  BUFX2 U19 ( .A(write), .Y(n2) );
  INVX1 U20 ( .A(N13), .Y(n167) );
  OR2X2 U21 ( .A(n96), .B(n58), .Y(n3) );
  AND2X2 U22 ( .A(n116), .B(n55), .Y(n4) );
  INVX1 U23 ( .A(n4), .Y(n5) );
  AND2X2 U24 ( .A(n113), .B(n55), .Y(n6) );
  INVX1 U25 ( .A(n6), .Y(n7) );
  AND2X2 U26 ( .A(n97), .B(n55), .Y(n8) );
  INVX1 U27 ( .A(n8), .Y(n9) );
  AND2X2 U28 ( .A(n100), .B(n55), .Y(n10) );
  INVX1 U29 ( .A(n10), .Y(n11) );
  AND2X2 U30 ( .A(n103), .B(n55), .Y(n12) );
  INVX1 U31 ( .A(n12), .Y(n13) );
  AND2X2 U32 ( .A(n106), .B(n55), .Y(n14) );
  INVX1 U33 ( .A(n14), .Y(n15) );
  AND2X2 U34 ( .A(n109), .B(n55), .Y(n16) );
  INVX1 U35 ( .A(n16), .Y(n17) );
  AND2X2 U36 ( .A(n115), .B(n55), .Y(n18) );
  INVX1 U37 ( .A(n18), .Y(n19) );
  AND2X2 U38 ( .A(n116), .B(n56), .Y(n20) );
  INVX1 U39 ( .A(n20), .Y(n21) );
  AND2X2 U40 ( .A(n113), .B(n56), .Y(n22) );
  INVX1 U41 ( .A(n22), .Y(n23) );
  AND2X2 U42 ( .A(n97), .B(n56), .Y(n24) );
  INVX1 U43 ( .A(n24), .Y(n25) );
  AND2X2 U44 ( .A(n100), .B(n56), .Y(n26) );
  INVX1 U45 ( .A(n26), .Y(n27) );
  AND2X2 U46 ( .A(n103), .B(n56), .Y(n28) );
  INVX1 U47 ( .A(n28), .Y(n29) );
  AND2X2 U48 ( .A(n106), .B(n56), .Y(n30) );
  INVX1 U49 ( .A(n30), .Y(n31) );
  AND2X2 U50 ( .A(n109), .B(n56), .Y(n32) );
  INVX1 U51 ( .A(n32), .Y(n33) );
  AND2X2 U52 ( .A(n115), .B(n56), .Y(n34) );
  INVX1 U53 ( .A(n34), .Y(n35) );
  INVX1 U54 ( .A(n36), .Y(n37) );
  INVX1 U55 ( .A(n38), .Y(n39) );
  INVX1 U56 ( .A(n40), .Y(n41) );
  INVX1 U57 ( .A(n42), .Y(n43) );
  INVX1 U58 ( .A(n44), .Y(n45) );
  INVX1 U59 ( .A(n46), .Y(n47) );
  INVX1 U60 ( .A(n48), .Y(n49) );
  INVX1 U61 ( .A(n50), .Y(n51) );
  OR2X2 U62 ( .A(\addr<5> ), .B(n3), .Y(n52) );
  INVX1 U63 ( .A(n52), .Y(n53) );
  INVX1 U64 ( .A(n52), .Y(n54) );
  AND2X2 U65 ( .A(\data_in<0> ), .B(n155), .Y(n55) );
  AND2X2 U66 ( .A(\data_in<0> ), .B(n153), .Y(n56) );
  AND2X2 U67 ( .A(\data_in<0> ), .B(n1), .Y(n57) );
  INVX1 U68 ( .A(n165), .Y(n164) );
  INVX1 U69 ( .A(n163), .Y(n162) );
  INVX1 U70 ( .A(n161), .Y(n160) );
  OR2X1 U71 ( .A(n59), .B(rst), .Y(n58) );
  OR2X1 U72 ( .A(\addr<6> ), .B(\addr<7> ), .Y(n59) );
  OR2X1 U73 ( .A(n162), .B(n164), .Y(n60) );
  INVX1 U74 ( .A(n60), .Y(n93) );
  INVX1 U75 ( .A(n186), .Y(n155) );
  INVX1 U76 ( .A(n209), .Y(n153) );
  AND2X1 U77 ( .A(n164), .B(n162), .Y(n94) );
  OR2X2 U78 ( .A(n3), .B(\addr<5> ), .Y(n95) );
  INVX1 U79 ( .A(write), .Y(n96) );
  INVX1 U80 ( .A(rst), .Y(n159) );
  INVX1 U81 ( .A(n99), .Y(n97) );
  INVX1 U82 ( .A(n97), .Y(n98) );
  BUFX2 U83 ( .A(n199), .Y(n99) );
  INVX1 U84 ( .A(n102), .Y(n100) );
  INVX1 U85 ( .A(n100), .Y(n101) );
  BUFX2 U86 ( .A(n201), .Y(n102) );
  INVX1 U87 ( .A(n105), .Y(n103) );
  INVX1 U88 ( .A(n103), .Y(n104) );
  BUFX2 U89 ( .A(n203), .Y(n105) );
  INVX1 U90 ( .A(n108), .Y(n106) );
  INVX1 U91 ( .A(n106), .Y(n107) );
  BUFX2 U92 ( .A(n205), .Y(n108) );
  INVX1 U94 ( .A(n111), .Y(n109) );
  INVX1 U95 ( .A(n109), .Y(n110) );
  BUFX2 U96 ( .A(n207), .Y(n111) );
  INVX1 U97 ( .A(n113), .Y(n112) );
  AND2X1 U98 ( .A(n161), .B(n94), .Y(n113) );
  INVX1 U99 ( .A(n115), .Y(n114) );
  AND2X1 U100 ( .A(n160), .B(n94), .Y(n116) );
  INVX1 U101 ( .A(n116), .Y(n117) );
  AND2X1 U102 ( .A(\data_in<0> ), .B(n157), .Y(n118) );
  INVX1 U103 ( .A(n118), .Y(n119) );
  MUX2X1 U104 ( .B(n121), .A(n122), .S(n151), .Y(n120) );
  MUX2X1 U105 ( .B(n124), .A(n125), .S(n151), .Y(n123) );
  MUX2X1 U106 ( .B(n127), .A(n128), .S(n151), .Y(n126) );
  MUX2X1 U107 ( .B(n130), .A(n131), .S(n151), .Y(n129) );
  MUX2X1 U108 ( .B(n133), .A(n134), .S(n166), .Y(n132) );
  MUX2X1 U109 ( .B(n136), .A(n137), .S(n151), .Y(n135) );
  MUX2X1 U110 ( .B(n139), .A(n140), .S(n151), .Y(n138) );
  MUX2X1 U111 ( .B(n142), .A(n143), .S(n151), .Y(n141) );
  MUX2X1 U112 ( .B(n145), .A(n146), .S(n151), .Y(n144) );
  MUX2X1 U113 ( .B(n148), .A(n149), .S(n166), .Y(n147) );
  MUX2X1 U114 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n152), .Y(n122) );
  MUX2X1 U115 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n152), .Y(n121) );
  MUX2X1 U116 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n152), .Y(n125) );
  MUX2X1 U117 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n152), .Y(n124) );
  MUX2X1 U118 ( .B(n123), .A(n120), .S(n164), .Y(n134) );
  MUX2X1 U119 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n152), .Y(n128) );
  MUX2X1 U120 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n152), .Y(n127) );
  MUX2X1 U121 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n152), .Y(n131) );
  MUX2X1 U122 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n152), .Y(n130) );
  MUX2X1 U123 ( .B(n129), .A(n126), .S(n164), .Y(n133) );
  MUX2X1 U124 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n152), .Y(n137) );
  MUX2X1 U125 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n152), .Y(n136) );
  MUX2X1 U126 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n152), .Y(n140) );
  MUX2X1 U127 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n152), .Y(n139) );
  MUX2X1 U128 ( .B(n138), .A(n135), .S(n164), .Y(n149) );
  MUX2X1 U129 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n152), .Y(n143) );
  MUX2X1 U130 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n152), .Y(n142) );
  MUX2X1 U131 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n152), .Y(n146) );
  MUX2X1 U132 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n152), .Y(n145) );
  MUX2X1 U133 ( .B(n144), .A(n141), .S(n164), .Y(n148) );
  MUX2X1 U134 ( .B(n147), .A(n132), .S(n168), .Y(n150) );
  INVX1 U135 ( .A(N12), .Y(n165) );
  INVX1 U136 ( .A(N11), .Y(n163) );
  INVX1 U137 ( .A(N10), .Y(n161) );
  NOR3X1 U138 ( .A(n169), .B(n167), .C(n95), .Y(n157) );
  INVX2 U139 ( .A(n157), .Y(n177) );
  INVX1 U140 ( .A(n169), .Y(n168) );
  INVX1 U141 ( .A(n167), .Y(n166) );
  OAI21X1 U142 ( .A(n177), .B(n117), .C(\mem<31><0> ), .Y(n170) );
  OAI21X1 U143 ( .A(n119), .B(n117), .C(n170), .Y(n61) );
  OAI21X1 U144 ( .A(n112), .B(n177), .C(\mem<30><0> ), .Y(n171) );
  OAI21X1 U145 ( .A(n112), .B(n119), .C(n171), .Y(n62) );
  NAND3X1 U146 ( .A(n160), .B(n164), .C(n163), .Y(n199) );
  OAI21X1 U147 ( .A(n98), .B(n177), .C(\mem<29><0> ), .Y(n172) );
  OAI21X1 U148 ( .A(n98), .B(n119), .C(n172), .Y(n63) );
  NAND3X1 U149 ( .A(n164), .B(n163), .C(n161), .Y(n201) );
  OAI21X1 U150 ( .A(n101), .B(n177), .C(\mem<28><0> ), .Y(n173) );
  OAI21X1 U151 ( .A(n101), .B(n119), .C(n173), .Y(n64) );
  NAND3X1 U152 ( .A(n160), .B(n162), .C(n165), .Y(n203) );
  OAI21X1 U153 ( .A(n104), .B(n177), .C(\mem<27><0> ), .Y(n174) );
  OAI21X1 U154 ( .A(n104), .B(n119), .C(n174), .Y(n65) );
  NAND3X1 U155 ( .A(n165), .B(n162), .C(n161), .Y(n205) );
  OAI21X1 U156 ( .A(n107), .B(n177), .C(\mem<26><0> ), .Y(n175) );
  OAI21X1 U157 ( .A(n107), .B(n119), .C(n175), .Y(n66) );
  NAND3X1 U158 ( .A(n160), .B(n165), .C(n163), .Y(n207) );
  OAI21X1 U159 ( .A(n110), .B(n177), .C(\mem<25><0> ), .Y(n176) );
  OAI21X1 U160 ( .A(n110), .B(n119), .C(n176), .Y(n67) );
  OAI21X1 U161 ( .A(n114), .B(n177), .C(\mem<24><0> ), .Y(n178) );
  OAI21X1 U162 ( .A(n114), .B(n119), .C(n178), .Y(n68) );
  NAND3X1 U163 ( .A(n54), .B(n168), .C(n167), .Y(n186) );
  OAI21X1 U164 ( .A(n156), .B(n117), .C(\mem<23><0> ), .Y(n179) );
  NAND2X1 U165 ( .A(n5), .B(n179), .Y(n69) );
  OAI21X1 U166 ( .A(n156), .B(n112), .C(\mem<22><0> ), .Y(n180) );
  NAND2X1 U167 ( .A(n7), .B(n180), .Y(n70) );
  OAI21X1 U168 ( .A(n156), .B(n98), .C(\mem<21><0> ), .Y(n181) );
  NAND2X1 U169 ( .A(n9), .B(n181), .Y(n71) );
  OAI21X1 U170 ( .A(n156), .B(n101), .C(\mem<20><0> ), .Y(n182) );
  NAND2X1 U171 ( .A(n11), .B(n182), .Y(n72) );
  OAI21X1 U172 ( .A(n156), .B(n104), .C(\mem<19><0> ), .Y(n183) );
  NAND2X1 U173 ( .A(n13), .B(n183), .Y(n73) );
  OAI21X1 U174 ( .A(n156), .B(n107), .C(\mem<18><0> ), .Y(n184) );
  NAND2X1 U175 ( .A(n15), .B(n184), .Y(n74) );
  OAI21X1 U176 ( .A(n156), .B(n110), .C(\mem<17><0> ), .Y(n185) );
  NAND2X1 U177 ( .A(n17), .B(n185), .Y(n75) );
  OAI21X1 U178 ( .A(n156), .B(n114), .C(\mem<16><0> ), .Y(n187) );
  NAND2X1 U179 ( .A(n19), .B(n187), .Y(n76) );
  OAI21X1 U180 ( .A(n195), .B(n117), .C(\mem<15><0> ), .Y(n188) );
  NAND2X1 U181 ( .A(n188), .B(n37), .Y(n77) );
  OAI21X1 U182 ( .A(n195), .B(n112), .C(\mem<14><0> ), .Y(n189) );
  NAND2X1 U183 ( .A(n39), .B(n189), .Y(n78) );
  OAI21X1 U184 ( .A(n195), .B(n98), .C(\mem<13><0> ), .Y(n190) );
  NAND2X1 U185 ( .A(n41), .B(n190), .Y(n79) );
  OAI21X1 U186 ( .A(n195), .B(n101), .C(\mem<12><0> ), .Y(n191) );
  NAND2X1 U187 ( .A(n43), .B(n191), .Y(n80) );
  OAI21X1 U188 ( .A(n195), .B(n104), .C(\mem<11><0> ), .Y(n192) );
  NAND2X1 U189 ( .A(n45), .B(n192), .Y(n81) );
  OAI21X1 U190 ( .A(n195), .B(n107), .C(\mem<10><0> ), .Y(n193) );
  NAND2X1 U191 ( .A(n47), .B(n193), .Y(n82) );
  OAI21X1 U192 ( .A(n195), .B(n110), .C(\mem<9><0> ), .Y(n194) );
  NAND2X1 U193 ( .A(n49), .B(n194), .Y(n83) );
  OAI21X1 U194 ( .A(n195), .B(n114), .C(\mem<8><0> ), .Y(n196) );
  NAND2X1 U195 ( .A(n51), .B(n196), .Y(n84) );
  NAND3X1 U196 ( .A(n53), .B(n167), .C(n169), .Y(n209) );
  OAI21X1 U197 ( .A(n154), .B(n117), .C(\mem<7><0> ), .Y(n197) );
  NAND2X1 U198 ( .A(n21), .B(n197), .Y(n85) );
  OAI21X1 U199 ( .A(n154), .B(n112), .C(\mem<6><0> ), .Y(n198) );
  NAND2X1 U200 ( .A(n23), .B(n198), .Y(n86) );
  OAI21X1 U201 ( .A(n154), .B(n98), .C(\mem<5><0> ), .Y(n200) );
  NAND2X1 U202 ( .A(n25), .B(n200), .Y(n87) );
  OAI21X1 U203 ( .A(n154), .B(n101), .C(\mem<4><0> ), .Y(n202) );
  NAND2X1 U204 ( .A(n27), .B(n202), .Y(n88) );
  OAI21X1 U205 ( .A(n154), .B(n104), .C(\mem<3><0> ), .Y(n204) );
  NAND2X1 U206 ( .A(n29), .B(n204), .Y(n89) );
  OAI21X1 U207 ( .A(n154), .B(n107), .C(\mem<2><0> ), .Y(n206) );
  NAND2X1 U208 ( .A(n31), .B(n206), .Y(n90) );
  OAI21X1 U209 ( .A(n154), .B(n110), .C(\mem<1><0> ), .Y(n208) );
  NAND2X1 U210 ( .A(n33), .B(n208), .Y(n91) );
  OAI21X1 U211 ( .A(n154), .B(n114), .C(\mem<0><0> ), .Y(n210) );
  NAND2X1 U212 ( .A(n35), .B(n210), .Y(n92) );
endmodule


module memv ( data_out, .addr({\addr<7> , \addr<6> , \addr<5> , \addr<4> , 
        \addr<3> , \addr<2> , \addr<1> , \addr<0> }), data_in, write, clk, rst, 
        createdump, .file_id({\file_id<4> , \file_id<3> , \file_id<2> , 
        \file_id<1> , \file_id<0> }) );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , data_in, write, clk, rst, createdump,
         \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> ;
  output data_out;
  wire   N18, N19, N20, N21, N22, N23, N24, N25, \mem<0> , \mem<1> , \mem<2> ,
         \mem<3> , \mem<4> , \mem<5> , \mem<6> , \mem<7> , \mem<8> , \mem<9> ,
         \mem<10> , \mem<11> , \mem<12> , \mem<13> , \mem<14> , \mem<15> ,
         \mem<16> , \mem<17> , \mem<18> , \mem<19> , \mem<20> , \mem<21> ,
         \mem<22> , \mem<23> , \mem<24> , \mem<25> , \mem<26> , \mem<27> ,
         \mem<28> , \mem<29> , \mem<30> , \mem<31> , \mem<32> , \mem<33> ,
         \mem<34> , \mem<35> , \mem<36> , \mem<37> , \mem<38> , \mem<39> ,
         \mem<40> , \mem<41> , \mem<42> , \mem<43> , \mem<44> , \mem<45> ,
         \mem<46> , \mem<47> , \mem<48> , \mem<49> , \mem<50> , \mem<51> ,
         \mem<52> , \mem<53> , \mem<54> , \mem<55> , \mem<56> , \mem<57> ,
         \mem<58> , \mem<59> , \mem<60> , \mem<61> , \mem<62> , \mem<63> ,
         \mem<64> , \mem<65> , \mem<66> , \mem<67> , \mem<68> , \mem<69> ,
         \mem<70> , \mem<71> , \mem<72> , \mem<73> , \mem<74> , \mem<75> ,
         \mem<76> , \mem<77> , \mem<78> , \mem<79> , \mem<80> , \mem<81> ,
         \mem<82> , \mem<83> , \mem<84> , \mem<85> , \mem<86> , \mem<87> ,
         \mem<88> , \mem<89> , \mem<90> , \mem<91> , \mem<92> , \mem<93> ,
         \mem<94> , \mem<95> , \mem<96> , \mem<97> , \mem<98> , \mem<99> ,
         \mem<100> , \mem<101> , \mem<102> , \mem<103> , \mem<104> ,
         \mem<105> , \mem<106> , \mem<107> , \mem<108> , \mem<109> ,
         \mem<110> , \mem<111> , \mem<112> , \mem<113> , \mem<114> ,
         \mem<115> , \mem<116> , \mem<117> , \mem<118> , \mem<119> ,
         \mem<120> , \mem<121> , \mem<122> , \mem<123> , \mem<124> ,
         \mem<125> , \mem<126> , \mem<127> , \mem<128> , \mem<129> ,
         \mem<130> , \mem<131> , \mem<132> , \mem<133> , \mem<134> ,
         \mem<135> , \mem<136> , \mem<137> , \mem<138> , \mem<139> ,
         \mem<140> , \mem<141> , \mem<142> , \mem<143> , \mem<144> ,
         \mem<145> , \mem<146> , \mem<147> , \mem<148> , \mem<149> ,
         \mem<150> , \mem<151> , \mem<152> , \mem<153> , \mem<154> ,
         \mem<155> , \mem<156> , \mem<157> , \mem<158> , \mem<159> ,
         \mem<160> , \mem<161> , \mem<162> , \mem<163> , \mem<164> ,
         \mem<165> , \mem<166> , \mem<167> , \mem<168> , \mem<169> ,
         \mem<170> , \mem<171> , \mem<172> , \mem<173> , \mem<174> ,
         \mem<175> , \mem<176> , \mem<177> , \mem<178> , \mem<179> ,
         \mem<180> , \mem<181> , \mem<182> , \mem<183> , \mem<184> ,
         \mem<185> , \mem<186> , \mem<187> , \mem<188> , \mem<189> ,
         \mem<190> , \mem<191> , \mem<192> , \mem<193> , \mem<194> ,
         \mem<195> , \mem<196> , \mem<197> , \mem<198> , \mem<199> ,
         \mem<200> , \mem<201> , \mem<202> , \mem<203> , \mem<204> ,
         \mem<205> , \mem<206> , \mem<207> , \mem<208> , \mem<209> ,
         \mem<210> , \mem<211> , \mem<212> , \mem<213> , \mem<214> ,
         \mem<215> , \mem<216> , \mem<217> , \mem<218> , \mem<219> ,
         \mem<220> , \mem<221> , \mem<222> , \mem<223> , \mem<224> ,
         \mem<225> , \mem<226> , \mem<227> , \mem<228> , \mem<229> ,
         \mem<230> , \mem<231> , \mem<232> , \mem<233> , \mem<234> ,
         \mem<235> , \mem<236> , \mem<237> , \mem<238> , \mem<239> ,
         \mem<240> , \mem<241> , \mem<242> , \mem<243> , \mem<244> ,
         \mem<245> , \mem<246> , \mem<247> , \mem<248> , \mem<249> ,
         \mem<250> , \mem<251> , \mem<252> , \mem<253> , \mem<254> ,
         \mem<255> , N28, n42, n46, n49, n52, n55, n58, n61, n64, n67, n70,
         n73, n76, n79, n82, n85, n88, n90, n91, n92, n94, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n113, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n132, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n151, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n170, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n188, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n206, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n224,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n243, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n261, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n279, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n297, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n316, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n334, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n352, n355, n356, n357, n358, n359, n361, n363, n364, n365,
         n366, n367, n368, n370, n371, n372, n373, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n43, n44, n45, n47, n48, n50, n51, n53, n54, n56, n57, n59, n60, n62,
         n63, n65, n66, n68, n69, n71, n72, n74, n75, n77, n78, n80, n81, n83,
         n84, n86, n87, n89, n93, n95, n112, n114, n130, n131, n133, n149,
         n150, n152, n169, n171, n187, n189, n205, n207, n223, n225, n241,
         n242, n244, n260, n262, n278, n280, n296, n298, n314, n315, n317,
         n333, n335, n351, n353, n354, n360, n362, n369, n374, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005;
  assign N18 = \addr<0> ;
  assign N19 = \addr<1> ;
  assign N20 = \addr<2> ;
  assign N21 = \addr<3> ;
  assign N22 = \addr<4> ;
  assign N23 = \addr<5> ;
  assign N24 = \addr<6> ;
  assign N25 = \addr<7> ;

  DFFPOSX1 \mem_reg<0>  ( .D(n633), .CLK(clk), .Q(\mem<0> ) );
  DFFPOSX1 \mem_reg<1>  ( .D(n632), .CLK(clk), .Q(\mem<1> ) );
  DFFPOSX1 \mem_reg<2>  ( .D(n631), .CLK(clk), .Q(\mem<2> ) );
  DFFPOSX1 \mem_reg<3>  ( .D(n630), .CLK(clk), .Q(\mem<3> ) );
  DFFPOSX1 \mem_reg<4>  ( .D(n629), .CLK(clk), .Q(\mem<4> ) );
  DFFPOSX1 \mem_reg<5>  ( .D(n628), .CLK(clk), .Q(\mem<5> ) );
  DFFPOSX1 \mem_reg<6>  ( .D(n627), .CLK(clk), .Q(\mem<6> ) );
  DFFPOSX1 \mem_reg<7>  ( .D(n626), .CLK(clk), .Q(\mem<7> ) );
  DFFPOSX1 \mem_reg<8>  ( .D(n625), .CLK(clk), .Q(\mem<8> ) );
  DFFPOSX1 \mem_reg<9>  ( .D(n624), .CLK(clk), .Q(\mem<9> ) );
  DFFPOSX1 \mem_reg<10>  ( .D(n623), .CLK(clk), .Q(\mem<10> ) );
  DFFPOSX1 \mem_reg<11>  ( .D(n622), .CLK(clk), .Q(\mem<11> ) );
  DFFPOSX1 \mem_reg<12>  ( .D(n621), .CLK(clk), .Q(\mem<12> ) );
  DFFPOSX1 \mem_reg<13>  ( .D(n620), .CLK(clk), .Q(\mem<13> ) );
  DFFPOSX1 \mem_reg<14>  ( .D(n619), .CLK(clk), .Q(\mem<14> ) );
  DFFPOSX1 \mem_reg<15>  ( .D(n618), .CLK(clk), .Q(\mem<15> ) );
  DFFPOSX1 \mem_reg<16>  ( .D(n617), .CLK(clk), .Q(\mem<16> ) );
  DFFPOSX1 \mem_reg<17>  ( .D(n616), .CLK(clk), .Q(\mem<17> ) );
  DFFPOSX1 \mem_reg<18>  ( .D(n615), .CLK(clk), .Q(\mem<18> ) );
  DFFPOSX1 \mem_reg<19>  ( .D(n614), .CLK(clk), .Q(\mem<19> ) );
  DFFPOSX1 \mem_reg<20>  ( .D(n613), .CLK(clk), .Q(\mem<20> ) );
  DFFPOSX1 \mem_reg<21>  ( .D(n612), .CLK(clk), .Q(\mem<21> ) );
  DFFPOSX1 \mem_reg<22>  ( .D(n611), .CLK(clk), .Q(\mem<22> ) );
  DFFPOSX1 \mem_reg<23>  ( .D(n610), .CLK(clk), .Q(\mem<23> ) );
  DFFPOSX1 \mem_reg<24>  ( .D(n609), .CLK(clk), .Q(\mem<24> ) );
  DFFPOSX1 \mem_reg<25>  ( .D(n608), .CLK(clk), .Q(\mem<25> ) );
  DFFPOSX1 \mem_reg<26>  ( .D(n607), .CLK(clk), .Q(\mem<26> ) );
  DFFPOSX1 \mem_reg<27>  ( .D(n606), .CLK(clk), .Q(\mem<27> ) );
  DFFPOSX1 \mem_reg<28>  ( .D(n605), .CLK(clk), .Q(\mem<28> ) );
  DFFPOSX1 \mem_reg<29>  ( .D(n604), .CLK(clk), .Q(\mem<29> ) );
  DFFPOSX1 \mem_reg<30>  ( .D(n603), .CLK(clk), .Q(\mem<30> ) );
  DFFPOSX1 \mem_reg<31>  ( .D(n602), .CLK(clk), .Q(\mem<31> ) );
  DFFPOSX1 \mem_reg<32>  ( .D(n601), .CLK(clk), .Q(\mem<32> ) );
  DFFPOSX1 \mem_reg<33>  ( .D(n600), .CLK(clk), .Q(\mem<33> ) );
  DFFPOSX1 \mem_reg<34>  ( .D(n599), .CLK(clk), .Q(\mem<34> ) );
  DFFPOSX1 \mem_reg<35>  ( .D(n598), .CLK(clk), .Q(\mem<35> ) );
  DFFPOSX1 \mem_reg<36>  ( .D(n597), .CLK(clk), .Q(\mem<36> ) );
  DFFPOSX1 \mem_reg<37>  ( .D(n596), .CLK(clk), .Q(\mem<37> ) );
  DFFPOSX1 \mem_reg<38>  ( .D(n595), .CLK(clk), .Q(\mem<38> ) );
  DFFPOSX1 \mem_reg<39>  ( .D(n594), .CLK(clk), .Q(\mem<39> ) );
  DFFPOSX1 \mem_reg<40>  ( .D(n593), .CLK(clk), .Q(\mem<40> ) );
  DFFPOSX1 \mem_reg<41>  ( .D(n592), .CLK(clk), .Q(\mem<41> ) );
  DFFPOSX1 \mem_reg<42>  ( .D(n591), .CLK(clk), .Q(\mem<42> ) );
  DFFPOSX1 \mem_reg<43>  ( .D(n590), .CLK(clk), .Q(\mem<43> ) );
  DFFPOSX1 \mem_reg<44>  ( .D(n589), .CLK(clk), .Q(\mem<44> ) );
  DFFPOSX1 \mem_reg<45>  ( .D(n588), .CLK(clk), .Q(\mem<45> ) );
  DFFPOSX1 \mem_reg<46>  ( .D(n587), .CLK(clk), .Q(\mem<46> ) );
  DFFPOSX1 \mem_reg<47>  ( .D(n586), .CLK(clk), .Q(\mem<47> ) );
  DFFPOSX1 \mem_reg<48>  ( .D(n585), .CLK(clk), .Q(\mem<48> ) );
  DFFPOSX1 \mem_reg<49>  ( .D(n584), .CLK(clk), .Q(\mem<49> ) );
  DFFPOSX1 \mem_reg<50>  ( .D(n583), .CLK(clk), .Q(\mem<50> ) );
  DFFPOSX1 \mem_reg<51>  ( .D(n582), .CLK(clk), .Q(\mem<51> ) );
  DFFPOSX1 \mem_reg<52>  ( .D(n581), .CLK(clk), .Q(\mem<52> ) );
  DFFPOSX1 \mem_reg<53>  ( .D(n580), .CLK(clk), .Q(\mem<53> ) );
  DFFPOSX1 \mem_reg<54>  ( .D(n579), .CLK(clk), .Q(\mem<54> ) );
  DFFPOSX1 \mem_reg<55>  ( .D(n578), .CLK(clk), .Q(\mem<55> ) );
  DFFPOSX1 \mem_reg<56>  ( .D(n577), .CLK(clk), .Q(\mem<56> ) );
  DFFPOSX1 \mem_reg<57>  ( .D(n576), .CLK(clk), .Q(\mem<57> ) );
  DFFPOSX1 \mem_reg<58>  ( .D(n575), .CLK(clk), .Q(\mem<58> ) );
  DFFPOSX1 \mem_reg<59>  ( .D(n574), .CLK(clk), .Q(\mem<59> ) );
  DFFPOSX1 \mem_reg<60>  ( .D(n573), .CLK(clk), .Q(\mem<60> ) );
  DFFPOSX1 \mem_reg<61>  ( .D(n572), .CLK(clk), .Q(\mem<61> ) );
  DFFPOSX1 \mem_reg<62>  ( .D(n571), .CLK(clk), .Q(\mem<62> ) );
  DFFPOSX1 \mem_reg<63>  ( .D(n570), .CLK(clk), .Q(\mem<63> ) );
  DFFPOSX1 \mem_reg<64>  ( .D(n569), .CLK(clk), .Q(\mem<64> ) );
  DFFPOSX1 \mem_reg<65>  ( .D(n568), .CLK(clk), .Q(\mem<65> ) );
  DFFPOSX1 \mem_reg<66>  ( .D(n567), .CLK(clk), .Q(\mem<66> ) );
  DFFPOSX1 \mem_reg<67>  ( .D(n566), .CLK(clk), .Q(\mem<67> ) );
  DFFPOSX1 \mem_reg<68>  ( .D(n565), .CLK(clk), .Q(\mem<68> ) );
  DFFPOSX1 \mem_reg<69>  ( .D(n564), .CLK(clk), .Q(\mem<69> ) );
  DFFPOSX1 \mem_reg<70>  ( .D(n563), .CLK(clk), .Q(\mem<70> ) );
  DFFPOSX1 \mem_reg<71>  ( .D(n562), .CLK(clk), .Q(\mem<71> ) );
  DFFPOSX1 \mem_reg<72>  ( .D(n561), .CLK(clk), .Q(\mem<72> ) );
  DFFPOSX1 \mem_reg<73>  ( .D(n560), .CLK(clk), .Q(\mem<73> ) );
  DFFPOSX1 \mem_reg<74>  ( .D(n559), .CLK(clk), .Q(\mem<74> ) );
  DFFPOSX1 \mem_reg<75>  ( .D(n558), .CLK(clk), .Q(\mem<75> ) );
  DFFPOSX1 \mem_reg<76>  ( .D(n557), .CLK(clk), .Q(\mem<76> ) );
  DFFPOSX1 \mem_reg<77>  ( .D(n556), .CLK(clk), .Q(\mem<77> ) );
  DFFPOSX1 \mem_reg<78>  ( .D(n555), .CLK(clk), .Q(\mem<78> ) );
  DFFPOSX1 \mem_reg<79>  ( .D(n554), .CLK(clk), .Q(\mem<79> ) );
  DFFPOSX1 \mem_reg<80>  ( .D(n553), .CLK(clk), .Q(\mem<80> ) );
  DFFPOSX1 \mem_reg<81>  ( .D(n552), .CLK(clk), .Q(\mem<81> ) );
  DFFPOSX1 \mem_reg<82>  ( .D(n551), .CLK(clk), .Q(\mem<82> ) );
  DFFPOSX1 \mem_reg<83>  ( .D(n550), .CLK(clk), .Q(\mem<83> ) );
  DFFPOSX1 \mem_reg<84>  ( .D(n549), .CLK(clk), .Q(\mem<84> ) );
  DFFPOSX1 \mem_reg<85>  ( .D(n548), .CLK(clk), .Q(\mem<85> ) );
  DFFPOSX1 \mem_reg<86>  ( .D(n547), .CLK(clk), .Q(\mem<86> ) );
  DFFPOSX1 \mem_reg<87>  ( .D(n546), .CLK(clk), .Q(\mem<87> ) );
  DFFPOSX1 \mem_reg<88>  ( .D(n545), .CLK(clk), .Q(\mem<88> ) );
  DFFPOSX1 \mem_reg<89>  ( .D(n544), .CLK(clk), .Q(\mem<89> ) );
  DFFPOSX1 \mem_reg<90>  ( .D(n543), .CLK(clk), .Q(\mem<90> ) );
  DFFPOSX1 \mem_reg<91>  ( .D(n542), .CLK(clk), .Q(\mem<91> ) );
  DFFPOSX1 \mem_reg<92>  ( .D(n541), .CLK(clk), .Q(\mem<92> ) );
  DFFPOSX1 \mem_reg<93>  ( .D(n540), .CLK(clk), .Q(\mem<93> ) );
  DFFPOSX1 \mem_reg<94>  ( .D(n539), .CLK(clk), .Q(\mem<94> ) );
  DFFPOSX1 \mem_reg<95>  ( .D(n538), .CLK(clk), .Q(\mem<95> ) );
  DFFPOSX1 \mem_reg<96>  ( .D(n537), .CLK(clk), .Q(\mem<96> ) );
  DFFPOSX1 \mem_reg<97>  ( .D(n536), .CLK(clk), .Q(\mem<97> ) );
  DFFPOSX1 \mem_reg<98>  ( .D(n535), .CLK(clk), .Q(\mem<98> ) );
  DFFPOSX1 \mem_reg<99>  ( .D(n534), .CLK(clk), .Q(\mem<99> ) );
  DFFPOSX1 \mem_reg<100>  ( .D(n533), .CLK(clk), .Q(\mem<100> ) );
  DFFPOSX1 \mem_reg<101>  ( .D(n532), .CLK(clk), .Q(\mem<101> ) );
  DFFPOSX1 \mem_reg<102>  ( .D(n531), .CLK(clk), .Q(\mem<102> ) );
  DFFPOSX1 \mem_reg<103>  ( .D(n530), .CLK(clk), .Q(\mem<103> ) );
  DFFPOSX1 \mem_reg<104>  ( .D(n529), .CLK(clk), .Q(\mem<104> ) );
  DFFPOSX1 \mem_reg<105>  ( .D(n528), .CLK(clk), .Q(\mem<105> ) );
  DFFPOSX1 \mem_reg<106>  ( .D(n527), .CLK(clk), .Q(\mem<106> ) );
  DFFPOSX1 \mem_reg<107>  ( .D(n526), .CLK(clk), .Q(\mem<107> ) );
  DFFPOSX1 \mem_reg<108>  ( .D(n525), .CLK(clk), .Q(\mem<108> ) );
  DFFPOSX1 \mem_reg<109>  ( .D(n524), .CLK(clk), .Q(\mem<109> ) );
  DFFPOSX1 \mem_reg<110>  ( .D(n523), .CLK(clk), .Q(\mem<110> ) );
  DFFPOSX1 \mem_reg<111>  ( .D(n522), .CLK(clk), .Q(\mem<111> ) );
  DFFPOSX1 \mem_reg<112>  ( .D(n521), .CLK(clk), .Q(\mem<112> ) );
  DFFPOSX1 \mem_reg<113>  ( .D(n520), .CLK(clk), .Q(\mem<113> ) );
  DFFPOSX1 \mem_reg<114>  ( .D(n519), .CLK(clk), .Q(\mem<114> ) );
  DFFPOSX1 \mem_reg<115>  ( .D(n518), .CLK(clk), .Q(\mem<115> ) );
  DFFPOSX1 \mem_reg<116>  ( .D(n517), .CLK(clk), .Q(\mem<116> ) );
  DFFPOSX1 \mem_reg<117>  ( .D(n516), .CLK(clk), .Q(\mem<117> ) );
  DFFPOSX1 \mem_reg<118>  ( .D(n515), .CLK(clk), .Q(\mem<118> ) );
  DFFPOSX1 \mem_reg<119>  ( .D(n514), .CLK(clk), .Q(\mem<119> ) );
  DFFPOSX1 \mem_reg<120>  ( .D(n513), .CLK(clk), .Q(\mem<120> ) );
  DFFPOSX1 \mem_reg<121>  ( .D(n512), .CLK(clk), .Q(\mem<121> ) );
  DFFPOSX1 \mem_reg<122>  ( .D(n511), .CLK(clk), .Q(\mem<122> ) );
  DFFPOSX1 \mem_reg<123>  ( .D(n510), .CLK(clk), .Q(\mem<123> ) );
  DFFPOSX1 \mem_reg<124>  ( .D(n509), .CLK(clk), .Q(\mem<124> ) );
  DFFPOSX1 \mem_reg<125>  ( .D(n508), .CLK(clk), .Q(\mem<125> ) );
  DFFPOSX1 \mem_reg<126>  ( .D(n507), .CLK(clk), .Q(\mem<126> ) );
  DFFPOSX1 \mem_reg<127>  ( .D(n506), .CLK(clk), .Q(\mem<127> ) );
  DFFPOSX1 \mem_reg<128>  ( .D(n505), .CLK(clk), .Q(\mem<128> ) );
  DFFPOSX1 \mem_reg<129>  ( .D(n504), .CLK(clk), .Q(\mem<129> ) );
  DFFPOSX1 \mem_reg<130>  ( .D(n503), .CLK(clk), .Q(\mem<130> ) );
  DFFPOSX1 \mem_reg<131>  ( .D(n502), .CLK(clk), .Q(\mem<131> ) );
  DFFPOSX1 \mem_reg<132>  ( .D(n501), .CLK(clk), .Q(\mem<132> ) );
  DFFPOSX1 \mem_reg<133>  ( .D(n500), .CLK(clk), .Q(\mem<133> ) );
  DFFPOSX1 \mem_reg<134>  ( .D(n499), .CLK(clk), .Q(\mem<134> ) );
  DFFPOSX1 \mem_reg<135>  ( .D(n498), .CLK(clk), .Q(\mem<135> ) );
  DFFPOSX1 \mem_reg<136>  ( .D(n497), .CLK(clk), .Q(\mem<136> ) );
  DFFPOSX1 \mem_reg<137>  ( .D(n496), .CLK(clk), .Q(\mem<137> ) );
  DFFPOSX1 \mem_reg<138>  ( .D(n495), .CLK(clk), .Q(\mem<138> ) );
  DFFPOSX1 \mem_reg<139>  ( .D(n494), .CLK(clk), .Q(\mem<139> ) );
  DFFPOSX1 \mem_reg<140>  ( .D(n493), .CLK(clk), .Q(\mem<140> ) );
  DFFPOSX1 \mem_reg<141>  ( .D(n492), .CLK(clk), .Q(\mem<141> ) );
  DFFPOSX1 \mem_reg<142>  ( .D(n491), .CLK(clk), .Q(\mem<142> ) );
  DFFPOSX1 \mem_reg<143>  ( .D(n490), .CLK(clk), .Q(\mem<143> ) );
  DFFPOSX1 \mem_reg<144>  ( .D(n489), .CLK(clk), .Q(\mem<144> ) );
  DFFPOSX1 \mem_reg<145>  ( .D(n488), .CLK(clk), .Q(\mem<145> ) );
  DFFPOSX1 \mem_reg<146>  ( .D(n487), .CLK(clk), .Q(\mem<146> ) );
  DFFPOSX1 \mem_reg<147>  ( .D(n486), .CLK(clk), .Q(\mem<147> ) );
  DFFPOSX1 \mem_reg<148>  ( .D(n485), .CLK(clk), .Q(\mem<148> ) );
  DFFPOSX1 \mem_reg<149>  ( .D(n484), .CLK(clk), .Q(\mem<149> ) );
  DFFPOSX1 \mem_reg<150>  ( .D(n483), .CLK(clk), .Q(\mem<150> ) );
  DFFPOSX1 \mem_reg<151>  ( .D(n482), .CLK(clk), .Q(\mem<151> ) );
  DFFPOSX1 \mem_reg<152>  ( .D(n481), .CLK(clk), .Q(\mem<152> ) );
  DFFPOSX1 \mem_reg<153>  ( .D(n480), .CLK(clk), .Q(\mem<153> ) );
  DFFPOSX1 \mem_reg<154>  ( .D(n479), .CLK(clk), .Q(\mem<154> ) );
  DFFPOSX1 \mem_reg<155>  ( .D(n478), .CLK(clk), .Q(\mem<155> ) );
  DFFPOSX1 \mem_reg<156>  ( .D(n477), .CLK(clk), .Q(\mem<156> ) );
  DFFPOSX1 \mem_reg<157>  ( .D(n476), .CLK(clk), .Q(\mem<157> ) );
  DFFPOSX1 \mem_reg<158>  ( .D(n475), .CLK(clk), .Q(\mem<158> ) );
  DFFPOSX1 \mem_reg<159>  ( .D(n474), .CLK(clk), .Q(\mem<159> ) );
  DFFPOSX1 \mem_reg<160>  ( .D(n473), .CLK(clk), .Q(\mem<160> ) );
  DFFPOSX1 \mem_reg<161>  ( .D(n472), .CLK(clk), .Q(\mem<161> ) );
  DFFPOSX1 \mem_reg<162>  ( .D(n471), .CLK(clk), .Q(\mem<162> ) );
  DFFPOSX1 \mem_reg<163>  ( .D(n470), .CLK(clk), .Q(\mem<163> ) );
  DFFPOSX1 \mem_reg<164>  ( .D(n469), .CLK(clk), .Q(\mem<164> ) );
  DFFPOSX1 \mem_reg<165>  ( .D(n468), .CLK(clk), .Q(\mem<165> ) );
  DFFPOSX1 \mem_reg<166>  ( .D(n467), .CLK(clk), .Q(\mem<166> ) );
  DFFPOSX1 \mem_reg<167>  ( .D(n466), .CLK(clk), .Q(\mem<167> ) );
  DFFPOSX1 \mem_reg<168>  ( .D(n465), .CLK(clk), .Q(\mem<168> ) );
  DFFPOSX1 \mem_reg<169>  ( .D(n464), .CLK(clk), .Q(\mem<169> ) );
  DFFPOSX1 \mem_reg<170>  ( .D(n463), .CLK(clk), .Q(\mem<170> ) );
  DFFPOSX1 \mem_reg<171>  ( .D(n462), .CLK(clk), .Q(\mem<171> ) );
  DFFPOSX1 \mem_reg<172>  ( .D(n461), .CLK(clk), .Q(\mem<172> ) );
  DFFPOSX1 \mem_reg<173>  ( .D(n460), .CLK(clk), .Q(\mem<173> ) );
  DFFPOSX1 \mem_reg<174>  ( .D(n459), .CLK(clk), .Q(\mem<174> ) );
  DFFPOSX1 \mem_reg<175>  ( .D(n458), .CLK(clk), .Q(\mem<175> ) );
  DFFPOSX1 \mem_reg<176>  ( .D(n457), .CLK(clk), .Q(\mem<176> ) );
  DFFPOSX1 \mem_reg<177>  ( .D(n456), .CLK(clk), .Q(\mem<177> ) );
  DFFPOSX1 \mem_reg<178>  ( .D(n455), .CLK(clk), .Q(\mem<178> ) );
  DFFPOSX1 \mem_reg<179>  ( .D(n454), .CLK(clk), .Q(\mem<179> ) );
  DFFPOSX1 \mem_reg<180>  ( .D(n453), .CLK(clk), .Q(\mem<180> ) );
  DFFPOSX1 \mem_reg<181>  ( .D(n452), .CLK(clk), .Q(\mem<181> ) );
  DFFPOSX1 \mem_reg<182>  ( .D(n451), .CLK(clk), .Q(\mem<182> ) );
  DFFPOSX1 \mem_reg<183>  ( .D(n450), .CLK(clk), .Q(\mem<183> ) );
  DFFPOSX1 \mem_reg<184>  ( .D(n449), .CLK(clk), .Q(\mem<184> ) );
  DFFPOSX1 \mem_reg<185>  ( .D(n448), .CLK(clk), .Q(\mem<185> ) );
  DFFPOSX1 \mem_reg<186>  ( .D(n447), .CLK(clk), .Q(\mem<186> ) );
  DFFPOSX1 \mem_reg<187>  ( .D(n446), .CLK(clk), .Q(\mem<187> ) );
  DFFPOSX1 \mem_reg<188>  ( .D(n445), .CLK(clk), .Q(\mem<188> ) );
  DFFPOSX1 \mem_reg<189>  ( .D(n444), .CLK(clk), .Q(\mem<189> ) );
  DFFPOSX1 \mem_reg<190>  ( .D(n443), .CLK(clk), .Q(\mem<190> ) );
  DFFPOSX1 \mem_reg<191>  ( .D(n442), .CLK(clk), .Q(\mem<191> ) );
  DFFPOSX1 \mem_reg<192>  ( .D(n441), .CLK(clk), .Q(\mem<192> ) );
  DFFPOSX1 \mem_reg<193>  ( .D(n440), .CLK(clk), .Q(\mem<193> ) );
  DFFPOSX1 \mem_reg<194>  ( .D(n439), .CLK(clk), .Q(\mem<194> ) );
  DFFPOSX1 \mem_reg<195>  ( .D(n438), .CLK(clk), .Q(\mem<195> ) );
  DFFPOSX1 \mem_reg<196>  ( .D(n437), .CLK(clk), .Q(\mem<196> ) );
  DFFPOSX1 \mem_reg<197>  ( .D(n436), .CLK(clk), .Q(\mem<197> ) );
  DFFPOSX1 \mem_reg<198>  ( .D(n435), .CLK(clk), .Q(\mem<198> ) );
  DFFPOSX1 \mem_reg<199>  ( .D(n434), .CLK(clk), .Q(\mem<199> ) );
  DFFPOSX1 \mem_reg<200>  ( .D(n433), .CLK(clk), .Q(\mem<200> ) );
  DFFPOSX1 \mem_reg<201>  ( .D(n432), .CLK(clk), .Q(\mem<201> ) );
  DFFPOSX1 \mem_reg<202>  ( .D(n431), .CLK(clk), .Q(\mem<202> ) );
  DFFPOSX1 \mem_reg<203>  ( .D(n430), .CLK(clk), .Q(\mem<203> ) );
  DFFPOSX1 \mem_reg<204>  ( .D(n429), .CLK(clk), .Q(\mem<204> ) );
  DFFPOSX1 \mem_reg<205>  ( .D(n428), .CLK(clk), .Q(\mem<205> ) );
  DFFPOSX1 \mem_reg<206>  ( .D(n427), .CLK(clk), .Q(\mem<206> ) );
  DFFPOSX1 \mem_reg<207>  ( .D(n426), .CLK(clk), .Q(\mem<207> ) );
  DFFPOSX1 \mem_reg<208>  ( .D(n425), .CLK(clk), .Q(\mem<208> ) );
  DFFPOSX1 \mem_reg<209>  ( .D(n424), .CLK(clk), .Q(\mem<209> ) );
  DFFPOSX1 \mem_reg<210>  ( .D(n423), .CLK(clk), .Q(\mem<210> ) );
  DFFPOSX1 \mem_reg<211>  ( .D(n422), .CLK(clk), .Q(\mem<211> ) );
  DFFPOSX1 \mem_reg<212>  ( .D(n421), .CLK(clk), .Q(\mem<212> ) );
  DFFPOSX1 \mem_reg<213>  ( .D(n420), .CLK(clk), .Q(\mem<213> ) );
  DFFPOSX1 \mem_reg<214>  ( .D(n419), .CLK(clk), .Q(\mem<214> ) );
  DFFPOSX1 \mem_reg<215>  ( .D(n418), .CLK(clk), .Q(\mem<215> ) );
  DFFPOSX1 \mem_reg<216>  ( .D(n417), .CLK(clk), .Q(\mem<216> ) );
  DFFPOSX1 \mem_reg<217>  ( .D(n416), .CLK(clk), .Q(\mem<217> ) );
  DFFPOSX1 \mem_reg<218>  ( .D(n415), .CLK(clk), .Q(\mem<218> ) );
  DFFPOSX1 \mem_reg<219>  ( .D(n414), .CLK(clk), .Q(\mem<219> ) );
  DFFPOSX1 \mem_reg<220>  ( .D(n413), .CLK(clk), .Q(\mem<220> ) );
  DFFPOSX1 \mem_reg<221>  ( .D(n412), .CLK(clk), .Q(\mem<221> ) );
  DFFPOSX1 \mem_reg<222>  ( .D(n411), .CLK(clk), .Q(\mem<222> ) );
  DFFPOSX1 \mem_reg<223>  ( .D(n410), .CLK(clk), .Q(\mem<223> ) );
  DFFPOSX1 \mem_reg<224>  ( .D(n409), .CLK(clk), .Q(\mem<224> ) );
  DFFPOSX1 \mem_reg<225>  ( .D(n408), .CLK(clk), .Q(\mem<225> ) );
  DFFPOSX1 \mem_reg<226>  ( .D(n407), .CLK(clk), .Q(\mem<226> ) );
  DFFPOSX1 \mem_reg<227>  ( .D(n406), .CLK(clk), .Q(\mem<227> ) );
  DFFPOSX1 \mem_reg<228>  ( .D(n405), .CLK(clk), .Q(\mem<228> ) );
  DFFPOSX1 \mem_reg<229>  ( .D(n404), .CLK(clk), .Q(\mem<229> ) );
  DFFPOSX1 \mem_reg<230>  ( .D(n403), .CLK(clk), .Q(\mem<230> ) );
  DFFPOSX1 \mem_reg<231>  ( .D(n402), .CLK(clk), .Q(\mem<231> ) );
  DFFPOSX1 \mem_reg<232>  ( .D(n401), .CLK(clk), .Q(\mem<232> ) );
  DFFPOSX1 \mem_reg<233>  ( .D(n400), .CLK(clk), .Q(\mem<233> ) );
  DFFPOSX1 \mem_reg<234>  ( .D(n399), .CLK(clk), .Q(\mem<234> ) );
  DFFPOSX1 \mem_reg<235>  ( .D(n398), .CLK(clk), .Q(\mem<235> ) );
  DFFPOSX1 \mem_reg<236>  ( .D(n397), .CLK(clk), .Q(\mem<236> ) );
  DFFPOSX1 \mem_reg<237>  ( .D(n396), .CLK(clk), .Q(\mem<237> ) );
  DFFPOSX1 \mem_reg<238>  ( .D(n395), .CLK(clk), .Q(\mem<238> ) );
  DFFPOSX1 \mem_reg<239>  ( .D(n394), .CLK(clk), .Q(\mem<239> ) );
  DFFPOSX1 \mem_reg<240>  ( .D(n393), .CLK(clk), .Q(\mem<240> ) );
  DFFPOSX1 \mem_reg<241>  ( .D(n392), .CLK(clk), .Q(\mem<241> ) );
  DFFPOSX1 \mem_reg<242>  ( .D(n391), .CLK(clk), .Q(\mem<242> ) );
  DFFPOSX1 \mem_reg<243>  ( .D(n390), .CLK(clk), .Q(\mem<243> ) );
  DFFPOSX1 \mem_reg<244>  ( .D(n389), .CLK(clk), .Q(\mem<244> ) );
  DFFPOSX1 \mem_reg<245>  ( .D(n388), .CLK(clk), .Q(\mem<245> ) );
  DFFPOSX1 \mem_reg<246>  ( .D(n387), .CLK(clk), .Q(\mem<246> ) );
  DFFPOSX1 \mem_reg<247>  ( .D(n386), .CLK(clk), .Q(\mem<247> ) );
  DFFPOSX1 \mem_reg<248>  ( .D(n385), .CLK(clk), .Q(\mem<248> ) );
  DFFPOSX1 \mem_reg<249>  ( .D(n384), .CLK(clk), .Q(\mem<249> ) );
  DFFPOSX1 \mem_reg<250>  ( .D(n383), .CLK(clk), .Q(\mem<250> ) );
  DFFPOSX1 \mem_reg<251>  ( .D(n382), .CLK(clk), .Q(\mem<251> ) );
  DFFPOSX1 \mem_reg<252>  ( .D(n381), .CLK(clk), .Q(\mem<252> ) );
  DFFPOSX1 \mem_reg<253>  ( .D(n380), .CLK(clk), .Q(\mem<253> ) );
  DFFPOSX1 \mem_reg<254>  ( .D(n379), .CLK(clk), .Q(\mem<254> ) );
  DFFPOSX1 \mem_reg<255>  ( .D(n378), .CLK(clk), .Q(\mem<255> ) );
  AND2X2 U6 ( .A(N21), .B(n905), .Y(n355) );
  AND2X2 U7 ( .A(N21), .B(n1000), .Y(n364) );
  OAI21X1 U49 ( .A(n81), .B(n992), .C(n42), .Y(n378) );
  OAI21X1 U50 ( .A(n32), .B(n990), .C(\mem<255> ), .Y(n42) );
  OAI21X1 U51 ( .A(n993), .B(n78), .C(n46), .Y(n379) );
  OAI21X1 U52 ( .A(n991), .B(n30), .C(\mem<254> ), .Y(n46) );
  OAI21X1 U53 ( .A(n993), .B(n942), .C(n49), .Y(n380) );
  OAI21X1 U54 ( .A(n991), .B(n28), .C(\mem<253> ), .Y(n49) );
  OAI21X1 U55 ( .A(n993), .B(n941), .C(n52), .Y(n381) );
  OAI21X1 U56 ( .A(n991), .B(n26), .C(\mem<252> ), .Y(n52) );
  OAI21X1 U57 ( .A(n993), .B(n75), .C(n55), .Y(n382) );
  OAI21X1 U58 ( .A(n991), .B(n24), .C(\mem<251> ), .Y(n55) );
  OAI21X1 U59 ( .A(n993), .B(n72), .C(n58), .Y(n383) );
  OAI21X1 U60 ( .A(n991), .B(n22), .C(\mem<250> ), .Y(n58) );
  OAI21X1 U61 ( .A(n993), .B(n69), .C(n61), .Y(n384) );
  OAI21X1 U62 ( .A(n991), .B(n20), .C(\mem<249> ), .Y(n61) );
  OAI21X1 U63 ( .A(n993), .B(n66), .C(n64), .Y(n385) );
  OAI21X1 U64 ( .A(n991), .B(n18), .C(\mem<248> ), .Y(n64) );
  OAI21X1 U65 ( .A(n993), .B(n940), .C(n67), .Y(n386) );
  OAI21X1 U66 ( .A(n991), .B(n16), .C(\mem<247> ), .Y(n67) );
  OAI21X1 U67 ( .A(n992), .B(n939), .C(n70), .Y(n387) );
  OAI21X1 U68 ( .A(n990), .B(n14), .C(\mem<246> ), .Y(n70) );
  OAI21X1 U69 ( .A(n992), .B(n938), .C(n73), .Y(n388) );
  OAI21X1 U70 ( .A(n990), .B(n12), .C(\mem<245> ), .Y(n73) );
  OAI21X1 U71 ( .A(n992), .B(n937), .C(n76), .Y(n389) );
  OAI21X1 U72 ( .A(n990), .B(n10), .C(\mem<244> ), .Y(n76) );
  OAI21X1 U73 ( .A(n992), .B(n936), .C(n79), .Y(n390) );
  OAI21X1 U74 ( .A(n990), .B(n8), .C(\mem<243> ), .Y(n79) );
  OAI21X1 U75 ( .A(n992), .B(n935), .C(n82), .Y(n391) );
  OAI21X1 U76 ( .A(n990), .B(n6), .C(\mem<242> ), .Y(n82) );
  OAI21X1 U77 ( .A(n992), .B(n934), .C(n85), .Y(n392) );
  OAI21X1 U78 ( .A(n990), .B(n4), .C(\mem<241> ), .Y(n85) );
  OAI21X1 U79 ( .A(n992), .B(n928), .C(n88), .Y(n393) );
  OAI21X1 U80 ( .A(n990), .B(n2), .C(\mem<240> ), .Y(n88) );
  OAI21X1 U83 ( .A(n81), .B(n989), .C(n94), .Y(n394) );
  OAI21X1 U84 ( .A(n32), .B(n987), .C(\mem<239> ), .Y(n94) );
  OAI21X1 U85 ( .A(n78), .B(n989), .C(n96), .Y(n395) );
  OAI21X1 U86 ( .A(n30), .B(n987), .C(\mem<238> ), .Y(n96) );
  OAI21X1 U87 ( .A(n942), .B(n989), .C(n97), .Y(n396) );
  OAI21X1 U88 ( .A(n28), .B(n987), .C(\mem<237> ), .Y(n97) );
  OAI21X1 U89 ( .A(n941), .B(n989), .C(n98), .Y(n397) );
  OAI21X1 U90 ( .A(n26), .B(n987), .C(\mem<236> ), .Y(n98) );
  OAI21X1 U91 ( .A(n75), .B(n989), .C(n99), .Y(n398) );
  OAI21X1 U92 ( .A(n24), .B(n987), .C(\mem<235> ), .Y(n99) );
  OAI21X1 U93 ( .A(n72), .B(n989), .C(n100), .Y(n399) );
  OAI21X1 U94 ( .A(n22), .B(n987), .C(\mem<234> ), .Y(n100) );
  OAI21X1 U95 ( .A(n69), .B(n989), .C(n101), .Y(n400) );
  OAI21X1 U96 ( .A(n20), .B(n987), .C(\mem<233> ), .Y(n101) );
  OAI21X1 U97 ( .A(n66), .B(n989), .C(n102), .Y(n401) );
  OAI21X1 U98 ( .A(n18), .B(n987), .C(\mem<232> ), .Y(n102) );
  OAI21X1 U99 ( .A(n940), .B(n988), .C(n103), .Y(n402) );
  OAI21X1 U100 ( .A(n16), .B(n986), .C(\mem<231> ), .Y(n103) );
  OAI21X1 U101 ( .A(n939), .B(n988), .C(n104), .Y(n403) );
  OAI21X1 U102 ( .A(n14), .B(n986), .C(\mem<230> ), .Y(n104) );
  OAI21X1 U103 ( .A(n938), .B(n988), .C(n105), .Y(n404) );
  OAI21X1 U104 ( .A(n12), .B(n986), .C(\mem<229> ), .Y(n105) );
  OAI21X1 U105 ( .A(n937), .B(n988), .C(n106), .Y(n405) );
  OAI21X1 U106 ( .A(n10), .B(n986), .C(\mem<228> ), .Y(n106) );
  OAI21X1 U107 ( .A(n936), .B(n988), .C(n107), .Y(n406) );
  OAI21X1 U108 ( .A(n8), .B(n986), .C(\mem<227> ), .Y(n107) );
  OAI21X1 U109 ( .A(n935), .B(n988), .C(n108), .Y(n407) );
  OAI21X1 U110 ( .A(n6), .B(n986), .C(\mem<226> ), .Y(n108) );
  OAI21X1 U111 ( .A(n934), .B(n988), .C(n109), .Y(n408) );
  OAI21X1 U112 ( .A(n4), .B(n986), .C(\mem<225> ), .Y(n109) );
  OAI21X1 U113 ( .A(n928), .B(n988), .C(n110), .Y(n409) );
  OAI21X1 U114 ( .A(n2), .B(n986), .C(\mem<224> ), .Y(n110) );
  OAI21X1 U117 ( .A(n81), .B(n985), .C(n113), .Y(n410) );
  OAI21X1 U118 ( .A(n32), .B(n983), .C(\mem<223> ), .Y(n113) );
  OAI21X1 U119 ( .A(n78), .B(n985), .C(n115), .Y(n411) );
  OAI21X1 U120 ( .A(n30), .B(n983), .C(\mem<222> ), .Y(n115) );
  OAI21X1 U121 ( .A(n942), .B(n985), .C(n116), .Y(n412) );
  OAI21X1 U122 ( .A(n28), .B(n983), .C(\mem<221> ), .Y(n116) );
  OAI21X1 U123 ( .A(n941), .B(n985), .C(n117), .Y(n413) );
  OAI21X1 U124 ( .A(n26), .B(n983), .C(\mem<220> ), .Y(n117) );
  OAI21X1 U125 ( .A(n75), .B(n985), .C(n118), .Y(n414) );
  OAI21X1 U126 ( .A(n24), .B(n983), .C(\mem<219> ), .Y(n118) );
  OAI21X1 U127 ( .A(n72), .B(n985), .C(n119), .Y(n415) );
  OAI21X1 U128 ( .A(n22), .B(n983), .C(\mem<218> ), .Y(n119) );
  OAI21X1 U129 ( .A(n69), .B(n985), .C(n120), .Y(n416) );
  OAI21X1 U130 ( .A(n20), .B(n983), .C(\mem<217> ), .Y(n120) );
  OAI21X1 U131 ( .A(n66), .B(n985), .C(n121), .Y(n417) );
  OAI21X1 U132 ( .A(n18), .B(n983), .C(\mem<216> ), .Y(n121) );
  OAI21X1 U133 ( .A(n940), .B(n984), .C(n122), .Y(n418) );
  OAI21X1 U134 ( .A(n16), .B(n983), .C(\mem<215> ), .Y(n122) );
  OAI21X1 U135 ( .A(n939), .B(n984), .C(n123), .Y(n419) );
  OAI21X1 U136 ( .A(n14), .B(n983), .C(\mem<214> ), .Y(n123) );
  OAI21X1 U137 ( .A(n938), .B(n984), .C(n124), .Y(n420) );
  OAI21X1 U138 ( .A(n12), .B(n983), .C(\mem<213> ), .Y(n124) );
  OAI21X1 U139 ( .A(n937), .B(n984), .C(n125), .Y(n421) );
  OAI21X1 U140 ( .A(n10), .B(n983), .C(\mem<212> ), .Y(n125) );
  OAI21X1 U141 ( .A(n936), .B(n984), .C(n126), .Y(n422) );
  OAI21X1 U142 ( .A(n8), .B(n983), .C(\mem<211> ), .Y(n126) );
  OAI21X1 U143 ( .A(n935), .B(n984), .C(n127), .Y(n423) );
  OAI21X1 U144 ( .A(n6), .B(n983), .C(\mem<210> ), .Y(n127) );
  OAI21X1 U145 ( .A(n934), .B(n984), .C(n128), .Y(n424) );
  OAI21X1 U146 ( .A(n4), .B(n983), .C(\mem<209> ), .Y(n128) );
  OAI21X1 U147 ( .A(n928), .B(n984), .C(n129), .Y(n425) );
  OAI21X1 U148 ( .A(n2), .B(n983), .C(\mem<208> ), .Y(n129) );
  OAI21X1 U151 ( .A(n81), .B(n982), .C(n132), .Y(n426) );
  OAI21X1 U152 ( .A(n32), .B(n980), .C(\mem<207> ), .Y(n132) );
  OAI21X1 U153 ( .A(n78), .B(n982), .C(n134), .Y(n427) );
  OAI21X1 U154 ( .A(n30), .B(n980), .C(\mem<206> ), .Y(n134) );
  OAI21X1 U155 ( .A(n942), .B(n982), .C(n135), .Y(n428) );
  OAI21X1 U156 ( .A(n28), .B(n980), .C(\mem<205> ), .Y(n135) );
  OAI21X1 U157 ( .A(n941), .B(n982), .C(n136), .Y(n429) );
  OAI21X1 U158 ( .A(n26), .B(n980), .C(\mem<204> ), .Y(n136) );
  OAI21X1 U159 ( .A(n75), .B(n982), .C(n137), .Y(n430) );
  OAI21X1 U160 ( .A(n24), .B(n980), .C(\mem<203> ), .Y(n137) );
  OAI21X1 U161 ( .A(n72), .B(n982), .C(n138), .Y(n431) );
  OAI21X1 U162 ( .A(n22), .B(n980), .C(\mem<202> ), .Y(n138) );
  OAI21X1 U163 ( .A(n69), .B(n982), .C(n139), .Y(n432) );
  OAI21X1 U164 ( .A(n20), .B(n980), .C(\mem<201> ), .Y(n139) );
  OAI21X1 U165 ( .A(n66), .B(n982), .C(n140), .Y(n433) );
  OAI21X1 U166 ( .A(n18), .B(n980), .C(\mem<200> ), .Y(n140) );
  OAI21X1 U167 ( .A(n940), .B(n981), .C(n141), .Y(n434) );
  OAI21X1 U168 ( .A(n16), .B(n980), .C(\mem<199> ), .Y(n141) );
  OAI21X1 U169 ( .A(n939), .B(n981), .C(n142), .Y(n435) );
  OAI21X1 U170 ( .A(n14), .B(n980), .C(\mem<198> ), .Y(n142) );
  OAI21X1 U171 ( .A(n938), .B(n981), .C(n143), .Y(n436) );
  OAI21X1 U172 ( .A(n12), .B(n980), .C(\mem<197> ), .Y(n143) );
  OAI21X1 U173 ( .A(n937), .B(n981), .C(n144), .Y(n437) );
  OAI21X1 U174 ( .A(n10), .B(n980), .C(\mem<196> ), .Y(n144) );
  OAI21X1 U175 ( .A(n936), .B(n981), .C(n145), .Y(n438) );
  OAI21X1 U176 ( .A(n8), .B(n980), .C(\mem<195> ), .Y(n145) );
  OAI21X1 U177 ( .A(n935), .B(n981), .C(n146), .Y(n439) );
  OAI21X1 U178 ( .A(n6), .B(n980), .C(\mem<194> ), .Y(n146) );
  OAI21X1 U179 ( .A(n934), .B(n981), .C(n147), .Y(n440) );
  OAI21X1 U180 ( .A(n4), .B(n980), .C(\mem<193> ), .Y(n147) );
  OAI21X1 U181 ( .A(n928), .B(n981), .C(n148), .Y(n441) );
  OAI21X1 U182 ( .A(n2), .B(n980), .C(\mem<192> ), .Y(n148) );
  OAI21X1 U185 ( .A(n81), .B(n979), .C(n151), .Y(n442) );
  OAI21X1 U186 ( .A(n32), .B(n977), .C(\mem<191> ), .Y(n151) );
  OAI21X1 U187 ( .A(n78), .B(n979), .C(n153), .Y(n443) );
  OAI21X1 U188 ( .A(n30), .B(n977), .C(\mem<190> ), .Y(n153) );
  OAI21X1 U189 ( .A(n942), .B(n979), .C(n154), .Y(n444) );
  OAI21X1 U190 ( .A(n28), .B(n977), .C(\mem<189> ), .Y(n154) );
  OAI21X1 U191 ( .A(n941), .B(n979), .C(n155), .Y(n445) );
  OAI21X1 U192 ( .A(n26), .B(n977), .C(\mem<188> ), .Y(n155) );
  OAI21X1 U193 ( .A(n75), .B(n979), .C(n156), .Y(n446) );
  OAI21X1 U194 ( .A(n24), .B(n977), .C(\mem<187> ), .Y(n156) );
  OAI21X1 U195 ( .A(n72), .B(n979), .C(n157), .Y(n447) );
  OAI21X1 U196 ( .A(n22), .B(n977), .C(\mem<186> ), .Y(n157) );
  OAI21X1 U197 ( .A(n69), .B(n979), .C(n158), .Y(n448) );
  OAI21X1 U198 ( .A(n20), .B(n977), .C(\mem<185> ), .Y(n158) );
  OAI21X1 U199 ( .A(n66), .B(n979), .C(n159), .Y(n449) );
  OAI21X1 U200 ( .A(n18), .B(n977), .C(\mem<184> ), .Y(n159) );
  OAI21X1 U201 ( .A(n940), .B(n978), .C(n160), .Y(n450) );
  OAI21X1 U202 ( .A(n16), .B(n976), .C(\mem<183> ), .Y(n160) );
  OAI21X1 U203 ( .A(n939), .B(n978), .C(n161), .Y(n451) );
  OAI21X1 U204 ( .A(n14), .B(n976), .C(\mem<182> ), .Y(n161) );
  OAI21X1 U205 ( .A(n938), .B(n978), .C(n162), .Y(n452) );
  OAI21X1 U206 ( .A(n12), .B(n976), .C(\mem<181> ), .Y(n162) );
  OAI21X1 U207 ( .A(n937), .B(n978), .C(n163), .Y(n453) );
  OAI21X1 U208 ( .A(n10), .B(n976), .C(\mem<180> ), .Y(n163) );
  OAI21X1 U209 ( .A(n936), .B(n978), .C(n164), .Y(n454) );
  OAI21X1 U210 ( .A(n8), .B(n976), .C(\mem<179> ), .Y(n164) );
  OAI21X1 U211 ( .A(n935), .B(n978), .C(n165), .Y(n455) );
  OAI21X1 U212 ( .A(n6), .B(n976), .C(\mem<178> ), .Y(n165) );
  OAI21X1 U213 ( .A(n934), .B(n978), .C(n166), .Y(n456) );
  OAI21X1 U214 ( .A(n4), .B(n976), .C(\mem<177> ), .Y(n166) );
  OAI21X1 U215 ( .A(n928), .B(n978), .C(n167), .Y(n457) );
  OAI21X1 U216 ( .A(n2), .B(n976), .C(\mem<176> ), .Y(n167) );
  OAI21X1 U219 ( .A(n81), .B(n975), .C(n170), .Y(n458) );
  OAI21X1 U220 ( .A(n32), .B(n973), .C(\mem<175> ), .Y(n170) );
  OAI21X1 U221 ( .A(n78), .B(n975), .C(n172), .Y(n459) );
  OAI21X1 U222 ( .A(n30), .B(n973), .C(\mem<174> ), .Y(n172) );
  OAI21X1 U223 ( .A(n942), .B(n975), .C(n173), .Y(n460) );
  OAI21X1 U224 ( .A(n28), .B(n973), .C(\mem<173> ), .Y(n173) );
  OAI21X1 U225 ( .A(n941), .B(n975), .C(n174), .Y(n461) );
  OAI21X1 U226 ( .A(n26), .B(n973), .C(\mem<172> ), .Y(n174) );
  OAI21X1 U227 ( .A(n75), .B(n975), .C(n175), .Y(n462) );
  OAI21X1 U228 ( .A(n24), .B(n973), .C(\mem<171> ), .Y(n175) );
  OAI21X1 U229 ( .A(n72), .B(n975), .C(n176), .Y(n463) );
  OAI21X1 U230 ( .A(n22), .B(n973), .C(\mem<170> ), .Y(n176) );
  OAI21X1 U231 ( .A(n69), .B(n975), .C(n177), .Y(n464) );
  OAI21X1 U232 ( .A(n20), .B(n973), .C(\mem<169> ), .Y(n177) );
  OAI21X1 U233 ( .A(n66), .B(n975), .C(n178), .Y(n465) );
  OAI21X1 U234 ( .A(n18), .B(n973), .C(\mem<168> ), .Y(n178) );
  OAI21X1 U235 ( .A(n940), .B(n974), .C(n179), .Y(n466) );
  OAI21X1 U236 ( .A(n16), .B(n972), .C(\mem<167> ), .Y(n179) );
  OAI21X1 U237 ( .A(n939), .B(n974), .C(n180), .Y(n467) );
  OAI21X1 U238 ( .A(n14), .B(n972), .C(\mem<166> ), .Y(n180) );
  OAI21X1 U239 ( .A(n938), .B(n974), .C(n181), .Y(n468) );
  OAI21X1 U240 ( .A(n12), .B(n972), .C(\mem<165> ), .Y(n181) );
  OAI21X1 U241 ( .A(n937), .B(n974), .C(n182), .Y(n469) );
  OAI21X1 U242 ( .A(n10), .B(n972), .C(\mem<164> ), .Y(n182) );
  OAI21X1 U243 ( .A(n936), .B(n974), .C(n183), .Y(n470) );
  OAI21X1 U244 ( .A(n8), .B(n972), .C(\mem<163> ), .Y(n183) );
  OAI21X1 U245 ( .A(n935), .B(n974), .C(n184), .Y(n471) );
  OAI21X1 U246 ( .A(n6), .B(n972), .C(\mem<162> ), .Y(n184) );
  OAI21X1 U247 ( .A(n934), .B(n974), .C(n185), .Y(n472) );
  OAI21X1 U248 ( .A(n4), .B(n972), .C(\mem<161> ), .Y(n185) );
  OAI21X1 U249 ( .A(n928), .B(n974), .C(n186), .Y(n473) );
  OAI21X1 U250 ( .A(n2), .B(n972), .C(\mem<160> ), .Y(n186) );
  OAI21X1 U253 ( .A(n81), .B(n971), .C(n188), .Y(n474) );
  OAI21X1 U254 ( .A(n32), .B(n969), .C(\mem<159> ), .Y(n188) );
  OAI21X1 U255 ( .A(n78), .B(n971), .C(n190), .Y(n475) );
  OAI21X1 U256 ( .A(n30), .B(n969), .C(\mem<158> ), .Y(n190) );
  OAI21X1 U257 ( .A(n942), .B(n971), .C(n191), .Y(n476) );
  OAI21X1 U258 ( .A(n28), .B(n969), .C(\mem<157> ), .Y(n191) );
  OAI21X1 U259 ( .A(n941), .B(n971), .C(n192), .Y(n477) );
  OAI21X1 U260 ( .A(n26), .B(n969), .C(\mem<156> ), .Y(n192) );
  OAI21X1 U261 ( .A(n75), .B(n971), .C(n193), .Y(n478) );
  OAI21X1 U262 ( .A(n24), .B(n969), .C(\mem<155> ), .Y(n193) );
  OAI21X1 U263 ( .A(n72), .B(n971), .C(n194), .Y(n479) );
  OAI21X1 U264 ( .A(n22), .B(n969), .C(\mem<154> ), .Y(n194) );
  OAI21X1 U265 ( .A(n69), .B(n971), .C(n195), .Y(n480) );
  OAI21X1 U266 ( .A(n20), .B(n969), .C(\mem<153> ), .Y(n195) );
  OAI21X1 U267 ( .A(n66), .B(n971), .C(n196), .Y(n481) );
  OAI21X1 U268 ( .A(n18), .B(n969), .C(\mem<152> ), .Y(n196) );
  OAI21X1 U269 ( .A(n940), .B(n970), .C(n197), .Y(n482) );
  OAI21X1 U270 ( .A(n16), .B(n968), .C(\mem<151> ), .Y(n197) );
  OAI21X1 U271 ( .A(n939), .B(n970), .C(n198), .Y(n483) );
  OAI21X1 U272 ( .A(n14), .B(n968), .C(\mem<150> ), .Y(n198) );
  OAI21X1 U273 ( .A(n938), .B(n970), .C(n199), .Y(n484) );
  OAI21X1 U274 ( .A(n12), .B(n968), .C(\mem<149> ), .Y(n199) );
  OAI21X1 U275 ( .A(n937), .B(n970), .C(n200), .Y(n485) );
  OAI21X1 U276 ( .A(n10), .B(n968), .C(\mem<148> ), .Y(n200) );
  OAI21X1 U277 ( .A(n936), .B(n970), .C(n201), .Y(n486) );
  OAI21X1 U278 ( .A(n8), .B(n968), .C(\mem<147> ), .Y(n201) );
  OAI21X1 U279 ( .A(n935), .B(n970), .C(n202), .Y(n487) );
  OAI21X1 U280 ( .A(n6), .B(n968), .C(\mem<146> ), .Y(n202) );
  OAI21X1 U281 ( .A(n934), .B(n970), .C(n203), .Y(n488) );
  OAI21X1 U282 ( .A(n4), .B(n968), .C(\mem<145> ), .Y(n203) );
  OAI21X1 U283 ( .A(n928), .B(n970), .C(n204), .Y(n489) );
  OAI21X1 U284 ( .A(n2), .B(n968), .C(\mem<144> ), .Y(n204) );
  OAI21X1 U287 ( .A(n81), .B(n967), .C(n206), .Y(n490) );
  OAI21X1 U288 ( .A(n32), .B(n965), .C(\mem<143> ), .Y(n206) );
  OAI21X1 U289 ( .A(n78), .B(n967), .C(n208), .Y(n491) );
  OAI21X1 U290 ( .A(n30), .B(n965), .C(\mem<142> ), .Y(n208) );
  OAI21X1 U291 ( .A(n942), .B(n967), .C(n209), .Y(n492) );
  OAI21X1 U292 ( .A(n28), .B(n965), .C(\mem<141> ), .Y(n209) );
  OAI21X1 U293 ( .A(n941), .B(n967), .C(n210), .Y(n493) );
  OAI21X1 U294 ( .A(n26), .B(n965), .C(\mem<140> ), .Y(n210) );
  OAI21X1 U295 ( .A(n75), .B(n967), .C(n211), .Y(n494) );
  OAI21X1 U296 ( .A(n24), .B(n965), .C(\mem<139> ), .Y(n211) );
  OAI21X1 U297 ( .A(n72), .B(n967), .C(n212), .Y(n495) );
  OAI21X1 U298 ( .A(n22), .B(n965), .C(\mem<138> ), .Y(n212) );
  OAI21X1 U299 ( .A(n69), .B(n967), .C(n213), .Y(n496) );
  OAI21X1 U300 ( .A(n20), .B(n965), .C(\mem<137> ), .Y(n213) );
  OAI21X1 U301 ( .A(n66), .B(n967), .C(n214), .Y(n497) );
  OAI21X1 U302 ( .A(n18), .B(n965), .C(\mem<136> ), .Y(n214) );
  OAI21X1 U303 ( .A(n940), .B(n966), .C(n215), .Y(n498) );
  OAI21X1 U304 ( .A(n16), .B(n964), .C(\mem<135> ), .Y(n215) );
  OAI21X1 U305 ( .A(n939), .B(n966), .C(n216), .Y(n499) );
  OAI21X1 U306 ( .A(n14), .B(n964), .C(\mem<134> ), .Y(n216) );
  OAI21X1 U307 ( .A(n938), .B(n966), .C(n217), .Y(n500) );
  OAI21X1 U308 ( .A(n12), .B(n964), .C(\mem<133> ), .Y(n217) );
  OAI21X1 U309 ( .A(n937), .B(n966), .C(n218), .Y(n501) );
  OAI21X1 U310 ( .A(n10), .B(n964), .C(\mem<132> ), .Y(n218) );
  OAI21X1 U311 ( .A(n936), .B(n966), .C(n219), .Y(n502) );
  OAI21X1 U312 ( .A(n8), .B(n964), .C(\mem<131> ), .Y(n219) );
  OAI21X1 U313 ( .A(n935), .B(n966), .C(n220), .Y(n503) );
  OAI21X1 U314 ( .A(n6), .B(n964), .C(\mem<130> ), .Y(n220) );
  OAI21X1 U315 ( .A(n934), .B(n966), .C(n221), .Y(n504) );
  OAI21X1 U316 ( .A(n4), .B(n964), .C(\mem<129> ), .Y(n221) );
  OAI21X1 U317 ( .A(n928), .B(n966), .C(n222), .Y(n505) );
  OAI21X1 U318 ( .A(n2), .B(n964), .C(\mem<128> ), .Y(n222) );
  OAI21X1 U321 ( .A(n81), .B(n963), .C(n224), .Y(n506) );
  OAI21X1 U322 ( .A(n32), .B(n961), .C(\mem<127> ), .Y(n224) );
  OAI21X1 U323 ( .A(n78), .B(n963), .C(n226), .Y(n507) );
  OAI21X1 U324 ( .A(n30), .B(n961), .C(\mem<126> ), .Y(n226) );
  OAI21X1 U325 ( .A(n942), .B(n963), .C(n227), .Y(n508) );
  OAI21X1 U326 ( .A(n28), .B(n961), .C(\mem<125> ), .Y(n227) );
  OAI21X1 U327 ( .A(n941), .B(n963), .C(n228), .Y(n509) );
  OAI21X1 U328 ( .A(n26), .B(n961), .C(\mem<124> ), .Y(n228) );
  OAI21X1 U329 ( .A(n75), .B(n963), .C(n229), .Y(n510) );
  OAI21X1 U330 ( .A(n24), .B(n961), .C(\mem<123> ), .Y(n229) );
  OAI21X1 U331 ( .A(n72), .B(n963), .C(n230), .Y(n511) );
  OAI21X1 U332 ( .A(n22), .B(n961), .C(\mem<122> ), .Y(n230) );
  OAI21X1 U333 ( .A(n69), .B(n963), .C(n231), .Y(n512) );
  OAI21X1 U334 ( .A(n20), .B(n961), .C(\mem<121> ), .Y(n231) );
  OAI21X1 U335 ( .A(n66), .B(n963), .C(n232), .Y(n513) );
  OAI21X1 U336 ( .A(n18), .B(n961), .C(\mem<120> ), .Y(n232) );
  OAI21X1 U337 ( .A(n940), .B(n962), .C(n233), .Y(n514) );
  OAI21X1 U338 ( .A(n16), .B(n961), .C(\mem<119> ), .Y(n233) );
  OAI21X1 U339 ( .A(n939), .B(n962), .C(n234), .Y(n515) );
  OAI21X1 U340 ( .A(n14), .B(n961), .C(\mem<118> ), .Y(n234) );
  OAI21X1 U341 ( .A(n938), .B(n962), .C(n235), .Y(n516) );
  OAI21X1 U342 ( .A(n12), .B(n961), .C(\mem<117> ), .Y(n235) );
  OAI21X1 U343 ( .A(n937), .B(n962), .C(n236), .Y(n517) );
  OAI21X1 U344 ( .A(n10), .B(n961), .C(\mem<116> ), .Y(n236) );
  OAI21X1 U345 ( .A(n936), .B(n962), .C(n237), .Y(n518) );
  OAI21X1 U346 ( .A(n8), .B(n961), .C(\mem<115> ), .Y(n237) );
  OAI21X1 U347 ( .A(n935), .B(n962), .C(n238), .Y(n519) );
  OAI21X1 U348 ( .A(n6), .B(n961), .C(\mem<114> ), .Y(n238) );
  OAI21X1 U349 ( .A(n934), .B(n962), .C(n239), .Y(n520) );
  OAI21X1 U350 ( .A(n4), .B(n961), .C(\mem<113> ), .Y(n239) );
  OAI21X1 U351 ( .A(n928), .B(n962), .C(n240), .Y(n521) );
  OAI21X1 U352 ( .A(n2), .B(n961), .C(\mem<112> ), .Y(n240) );
  OAI21X1 U355 ( .A(n81), .B(n960), .C(n243), .Y(n522) );
  OAI21X1 U356 ( .A(n32), .B(n958), .C(\mem<111> ), .Y(n243) );
  OAI21X1 U357 ( .A(n78), .B(n960), .C(n245), .Y(n523) );
  OAI21X1 U358 ( .A(n30), .B(n958), .C(\mem<110> ), .Y(n245) );
  OAI21X1 U359 ( .A(n942), .B(n960), .C(n246), .Y(n524) );
  OAI21X1 U360 ( .A(n28), .B(n958), .C(\mem<109> ), .Y(n246) );
  OAI21X1 U361 ( .A(n941), .B(n960), .C(n247), .Y(n525) );
  OAI21X1 U362 ( .A(n26), .B(n958), .C(\mem<108> ), .Y(n247) );
  OAI21X1 U363 ( .A(n75), .B(n960), .C(n248), .Y(n526) );
  OAI21X1 U364 ( .A(n24), .B(n958), .C(\mem<107> ), .Y(n248) );
  OAI21X1 U365 ( .A(n72), .B(n960), .C(n249), .Y(n527) );
  OAI21X1 U366 ( .A(n22), .B(n958), .C(\mem<106> ), .Y(n249) );
  OAI21X1 U367 ( .A(n69), .B(n960), .C(n250), .Y(n528) );
  OAI21X1 U368 ( .A(n20), .B(n958), .C(\mem<105> ), .Y(n250) );
  OAI21X1 U369 ( .A(n66), .B(n960), .C(n251), .Y(n529) );
  OAI21X1 U370 ( .A(n18), .B(n958), .C(\mem<104> ), .Y(n251) );
  OAI21X1 U371 ( .A(n940), .B(n959), .C(n252), .Y(n530) );
  OAI21X1 U372 ( .A(n16), .B(n958), .C(\mem<103> ), .Y(n252) );
  OAI21X1 U373 ( .A(n939), .B(n959), .C(n253), .Y(n531) );
  OAI21X1 U374 ( .A(n14), .B(n958), .C(\mem<102> ), .Y(n253) );
  OAI21X1 U375 ( .A(n938), .B(n959), .C(n254), .Y(n532) );
  OAI21X1 U376 ( .A(n12), .B(n958), .C(\mem<101> ), .Y(n254) );
  OAI21X1 U377 ( .A(n937), .B(n959), .C(n255), .Y(n533) );
  OAI21X1 U378 ( .A(n10), .B(n958), .C(\mem<100> ), .Y(n255) );
  OAI21X1 U379 ( .A(n936), .B(n959), .C(n256), .Y(n534) );
  OAI21X1 U380 ( .A(n8), .B(n958), .C(\mem<99> ), .Y(n256) );
  OAI21X1 U381 ( .A(n935), .B(n959), .C(n257), .Y(n535) );
  OAI21X1 U382 ( .A(n6), .B(n958), .C(\mem<98> ), .Y(n257) );
  OAI21X1 U383 ( .A(n934), .B(n959), .C(n258), .Y(n536) );
  OAI21X1 U384 ( .A(n4), .B(n958), .C(\mem<97> ), .Y(n258) );
  OAI21X1 U385 ( .A(n928), .B(n959), .C(n259), .Y(n537) );
  OAI21X1 U386 ( .A(n2), .B(n958), .C(\mem<96> ), .Y(n259) );
  OAI21X1 U389 ( .A(n81), .B(n957), .C(n261), .Y(n538) );
  OAI21X1 U390 ( .A(n32), .B(n955), .C(\mem<95> ), .Y(n261) );
  OAI21X1 U391 ( .A(n78), .B(n957), .C(n263), .Y(n539) );
  OAI21X1 U392 ( .A(n30), .B(n955), .C(\mem<94> ), .Y(n263) );
  OAI21X1 U393 ( .A(n942), .B(n957), .C(n264), .Y(n540) );
  OAI21X1 U394 ( .A(n28), .B(n955), .C(\mem<93> ), .Y(n264) );
  OAI21X1 U395 ( .A(n941), .B(n957), .C(n265), .Y(n541) );
  OAI21X1 U396 ( .A(n26), .B(n955), .C(\mem<92> ), .Y(n265) );
  OAI21X1 U397 ( .A(n75), .B(n957), .C(n266), .Y(n542) );
  OAI21X1 U398 ( .A(n24), .B(n955), .C(\mem<91> ), .Y(n266) );
  OAI21X1 U399 ( .A(n72), .B(n957), .C(n267), .Y(n543) );
  OAI21X1 U400 ( .A(n22), .B(n955), .C(\mem<90> ), .Y(n267) );
  OAI21X1 U401 ( .A(n69), .B(n957), .C(n268), .Y(n544) );
  OAI21X1 U402 ( .A(n20), .B(n955), .C(\mem<89> ), .Y(n268) );
  OAI21X1 U403 ( .A(n66), .B(n957), .C(n269), .Y(n545) );
  OAI21X1 U404 ( .A(n18), .B(n955), .C(\mem<88> ), .Y(n269) );
  OAI21X1 U405 ( .A(n940), .B(n956), .C(n270), .Y(n546) );
  OAI21X1 U406 ( .A(n16), .B(n955), .C(\mem<87> ), .Y(n270) );
  OAI21X1 U407 ( .A(n939), .B(n956), .C(n271), .Y(n547) );
  OAI21X1 U408 ( .A(n14), .B(n955), .C(\mem<86> ), .Y(n271) );
  OAI21X1 U409 ( .A(n938), .B(n956), .C(n272), .Y(n548) );
  OAI21X1 U410 ( .A(n12), .B(n955), .C(\mem<85> ), .Y(n272) );
  OAI21X1 U411 ( .A(n937), .B(n956), .C(n273), .Y(n549) );
  OAI21X1 U412 ( .A(n10), .B(n955), .C(\mem<84> ), .Y(n273) );
  OAI21X1 U413 ( .A(n936), .B(n956), .C(n274), .Y(n550) );
  OAI21X1 U414 ( .A(n8), .B(n955), .C(\mem<83> ), .Y(n274) );
  OAI21X1 U415 ( .A(n935), .B(n956), .C(n275), .Y(n551) );
  OAI21X1 U416 ( .A(n6), .B(n955), .C(\mem<82> ), .Y(n275) );
  OAI21X1 U417 ( .A(n934), .B(n956), .C(n276), .Y(n552) );
  OAI21X1 U418 ( .A(n4), .B(n955), .C(\mem<81> ), .Y(n276) );
  OAI21X1 U419 ( .A(n928), .B(n956), .C(n277), .Y(n553) );
  OAI21X1 U420 ( .A(n2), .B(n955), .C(\mem<80> ), .Y(n277) );
  OAI21X1 U423 ( .A(n81), .B(n954), .C(n279), .Y(n554) );
  OAI21X1 U424 ( .A(n32), .B(n952), .C(\mem<79> ), .Y(n279) );
  OAI21X1 U425 ( .A(n78), .B(n954), .C(n281), .Y(n555) );
  OAI21X1 U426 ( .A(n30), .B(n952), .C(\mem<78> ), .Y(n281) );
  OAI21X1 U427 ( .A(n942), .B(n954), .C(n282), .Y(n556) );
  OAI21X1 U428 ( .A(n28), .B(n952), .C(\mem<77> ), .Y(n282) );
  OAI21X1 U429 ( .A(n941), .B(n954), .C(n283), .Y(n557) );
  OAI21X1 U430 ( .A(n26), .B(n952), .C(\mem<76> ), .Y(n283) );
  OAI21X1 U431 ( .A(n75), .B(n954), .C(n284), .Y(n558) );
  OAI21X1 U432 ( .A(n24), .B(n952), .C(\mem<75> ), .Y(n284) );
  OAI21X1 U433 ( .A(n72), .B(n954), .C(n285), .Y(n559) );
  OAI21X1 U434 ( .A(n22), .B(n952), .C(\mem<74> ), .Y(n285) );
  OAI21X1 U435 ( .A(n69), .B(n954), .C(n286), .Y(n560) );
  OAI21X1 U436 ( .A(n20), .B(n952), .C(\mem<73> ), .Y(n286) );
  OAI21X1 U437 ( .A(n66), .B(n954), .C(n287), .Y(n561) );
  OAI21X1 U438 ( .A(n18), .B(n952), .C(\mem<72> ), .Y(n287) );
  OAI21X1 U439 ( .A(n940), .B(n953), .C(n288), .Y(n562) );
  OAI21X1 U440 ( .A(n16), .B(n952), .C(\mem<71> ), .Y(n288) );
  OAI21X1 U441 ( .A(n939), .B(n953), .C(n289), .Y(n563) );
  OAI21X1 U442 ( .A(n14), .B(n952), .C(\mem<70> ), .Y(n289) );
  OAI21X1 U443 ( .A(n938), .B(n953), .C(n290), .Y(n564) );
  OAI21X1 U444 ( .A(n12), .B(n952), .C(\mem<69> ), .Y(n290) );
  OAI21X1 U445 ( .A(n937), .B(n953), .C(n291), .Y(n565) );
  OAI21X1 U446 ( .A(n10), .B(n952), .C(\mem<68> ), .Y(n291) );
  OAI21X1 U447 ( .A(n936), .B(n953), .C(n292), .Y(n566) );
  OAI21X1 U448 ( .A(n8), .B(n952), .C(\mem<67> ), .Y(n292) );
  OAI21X1 U449 ( .A(n935), .B(n953), .C(n293), .Y(n567) );
  OAI21X1 U450 ( .A(n6), .B(n952), .C(\mem<66> ), .Y(n293) );
  OAI21X1 U451 ( .A(n934), .B(n953), .C(n294), .Y(n568) );
  OAI21X1 U452 ( .A(n4), .B(n952), .C(\mem<65> ), .Y(n294) );
  OAI21X1 U453 ( .A(n928), .B(n953), .C(n295), .Y(n569) );
  OAI21X1 U454 ( .A(n2), .B(n952), .C(\mem<64> ), .Y(n295) );
  OAI21X1 U458 ( .A(n81), .B(n951), .C(n297), .Y(n570) );
  OAI21X1 U459 ( .A(n32), .B(n949), .C(\mem<63> ), .Y(n297) );
  OAI21X1 U460 ( .A(n78), .B(n951), .C(n299), .Y(n571) );
  OAI21X1 U461 ( .A(n30), .B(n949), .C(\mem<62> ), .Y(n299) );
  OAI21X1 U462 ( .A(n942), .B(n951), .C(n300), .Y(n572) );
  OAI21X1 U463 ( .A(n28), .B(n949), .C(\mem<61> ), .Y(n300) );
  OAI21X1 U464 ( .A(n941), .B(n951), .C(n301), .Y(n573) );
  OAI21X1 U465 ( .A(n26), .B(n949), .C(\mem<60> ), .Y(n301) );
  OAI21X1 U466 ( .A(n75), .B(n951), .C(n302), .Y(n574) );
  OAI21X1 U467 ( .A(n24), .B(n949), .C(\mem<59> ), .Y(n302) );
  OAI21X1 U468 ( .A(n72), .B(n951), .C(n303), .Y(n575) );
  OAI21X1 U469 ( .A(n22), .B(n949), .C(\mem<58> ), .Y(n303) );
  OAI21X1 U470 ( .A(n69), .B(n951), .C(n304), .Y(n576) );
  OAI21X1 U471 ( .A(n20), .B(n949), .C(\mem<57> ), .Y(n304) );
  OAI21X1 U472 ( .A(n66), .B(n951), .C(n305), .Y(n577) );
  OAI21X1 U473 ( .A(n18), .B(n949), .C(\mem<56> ), .Y(n305) );
  OAI21X1 U474 ( .A(n940), .B(n950), .C(n306), .Y(n578) );
  OAI21X1 U475 ( .A(n16), .B(n949), .C(\mem<55> ), .Y(n306) );
  OAI21X1 U476 ( .A(n939), .B(n950), .C(n307), .Y(n579) );
  OAI21X1 U477 ( .A(n14), .B(n949), .C(\mem<54> ), .Y(n307) );
  OAI21X1 U478 ( .A(n938), .B(n950), .C(n308), .Y(n580) );
  OAI21X1 U479 ( .A(n12), .B(n949), .C(\mem<53> ), .Y(n308) );
  OAI21X1 U480 ( .A(n937), .B(n950), .C(n309), .Y(n581) );
  OAI21X1 U481 ( .A(n10), .B(n949), .C(\mem<52> ), .Y(n309) );
  OAI21X1 U482 ( .A(n936), .B(n950), .C(n310), .Y(n582) );
  OAI21X1 U483 ( .A(n8), .B(n949), .C(\mem<51> ), .Y(n310) );
  OAI21X1 U484 ( .A(n935), .B(n950), .C(n311), .Y(n583) );
  OAI21X1 U485 ( .A(n6), .B(n949), .C(\mem<50> ), .Y(n311) );
  OAI21X1 U486 ( .A(n934), .B(n950), .C(n312), .Y(n584) );
  OAI21X1 U487 ( .A(n4), .B(n949), .C(\mem<49> ), .Y(n312) );
  OAI21X1 U488 ( .A(n928), .B(n950), .C(n313), .Y(n585) );
  OAI21X1 U489 ( .A(n2), .B(n949), .C(\mem<48> ), .Y(n313) );
  OAI21X1 U492 ( .A(n81), .B(n948), .C(n316), .Y(n586) );
  OAI21X1 U493 ( .A(n32), .B(n946), .C(\mem<47> ), .Y(n316) );
  OAI21X1 U494 ( .A(n78), .B(n948), .C(n318), .Y(n587) );
  OAI21X1 U495 ( .A(n30), .B(n946), .C(\mem<46> ), .Y(n318) );
  OAI21X1 U496 ( .A(n942), .B(n948), .C(n319), .Y(n588) );
  OAI21X1 U497 ( .A(n28), .B(n946), .C(\mem<45> ), .Y(n319) );
  OAI21X1 U498 ( .A(n941), .B(n948), .C(n320), .Y(n589) );
  OAI21X1 U499 ( .A(n26), .B(n946), .C(\mem<44> ), .Y(n320) );
  OAI21X1 U500 ( .A(n75), .B(n948), .C(n321), .Y(n590) );
  OAI21X1 U501 ( .A(n24), .B(n946), .C(\mem<43> ), .Y(n321) );
  OAI21X1 U502 ( .A(n72), .B(n948), .C(n322), .Y(n591) );
  OAI21X1 U503 ( .A(n22), .B(n946), .C(\mem<42> ), .Y(n322) );
  OAI21X1 U504 ( .A(n69), .B(n948), .C(n323), .Y(n592) );
  OAI21X1 U505 ( .A(n20), .B(n946), .C(\mem<41> ), .Y(n323) );
  OAI21X1 U506 ( .A(n66), .B(n948), .C(n324), .Y(n593) );
  OAI21X1 U507 ( .A(n18), .B(n946), .C(\mem<40> ), .Y(n324) );
  OAI21X1 U508 ( .A(n940), .B(n947), .C(n325), .Y(n594) );
  OAI21X1 U509 ( .A(n16), .B(n946), .C(\mem<39> ), .Y(n325) );
  OAI21X1 U510 ( .A(n939), .B(n947), .C(n326), .Y(n595) );
  OAI21X1 U511 ( .A(n14), .B(n946), .C(\mem<38> ), .Y(n326) );
  OAI21X1 U512 ( .A(n938), .B(n947), .C(n327), .Y(n596) );
  OAI21X1 U513 ( .A(n12), .B(n946), .C(\mem<37> ), .Y(n327) );
  OAI21X1 U514 ( .A(n937), .B(n947), .C(n328), .Y(n597) );
  OAI21X1 U515 ( .A(n10), .B(n946), .C(\mem<36> ), .Y(n328) );
  OAI21X1 U516 ( .A(n936), .B(n947), .C(n329), .Y(n598) );
  OAI21X1 U517 ( .A(n8), .B(n946), .C(\mem<35> ), .Y(n329) );
  OAI21X1 U518 ( .A(n935), .B(n947), .C(n330), .Y(n599) );
  OAI21X1 U519 ( .A(n6), .B(n946), .C(\mem<34> ), .Y(n330) );
  OAI21X1 U520 ( .A(n934), .B(n947), .C(n331), .Y(n600) );
  OAI21X1 U521 ( .A(n4), .B(n946), .C(\mem<33> ), .Y(n331) );
  OAI21X1 U522 ( .A(n928), .B(n947), .C(n332), .Y(n601) );
  OAI21X1 U523 ( .A(n2), .B(n946), .C(\mem<32> ), .Y(n332) );
  OAI21X1 U526 ( .A(n81), .B(n945), .C(n334), .Y(n602) );
  OAI21X1 U527 ( .A(n32), .B(n943), .C(\mem<31> ), .Y(n334) );
  OAI21X1 U528 ( .A(n78), .B(n945), .C(n336), .Y(n603) );
  OAI21X1 U529 ( .A(n30), .B(n943), .C(\mem<30> ), .Y(n336) );
  OAI21X1 U530 ( .A(n942), .B(n945), .C(n337), .Y(n604) );
  OAI21X1 U531 ( .A(n28), .B(n943), .C(\mem<29> ), .Y(n337) );
  OAI21X1 U532 ( .A(n941), .B(n945), .C(n338), .Y(n605) );
  OAI21X1 U533 ( .A(n26), .B(n943), .C(\mem<28> ), .Y(n338) );
  OAI21X1 U534 ( .A(n75), .B(n945), .C(n339), .Y(n606) );
  OAI21X1 U535 ( .A(n24), .B(n943), .C(\mem<27> ), .Y(n339) );
  OAI21X1 U536 ( .A(n72), .B(n945), .C(n340), .Y(n607) );
  OAI21X1 U537 ( .A(n22), .B(n943), .C(\mem<26> ), .Y(n340) );
  OAI21X1 U538 ( .A(n69), .B(n945), .C(n341), .Y(n608) );
  OAI21X1 U539 ( .A(n20), .B(n943), .C(\mem<25> ), .Y(n341) );
  OAI21X1 U540 ( .A(n66), .B(n945), .C(n342), .Y(n609) );
  OAI21X1 U541 ( .A(n18), .B(n943), .C(\mem<24> ), .Y(n342) );
  OAI21X1 U542 ( .A(n940), .B(n944), .C(n343), .Y(n610) );
  OAI21X1 U543 ( .A(n16), .B(n943), .C(\mem<23> ), .Y(n343) );
  OAI21X1 U544 ( .A(n939), .B(n944), .C(n344), .Y(n611) );
  OAI21X1 U545 ( .A(n14), .B(n943), .C(\mem<22> ), .Y(n344) );
  OAI21X1 U546 ( .A(n938), .B(n944), .C(n345), .Y(n612) );
  OAI21X1 U547 ( .A(n12), .B(n943), .C(\mem<21> ), .Y(n345) );
  OAI21X1 U548 ( .A(n937), .B(n944), .C(n346), .Y(n613) );
  OAI21X1 U549 ( .A(n10), .B(n943), .C(\mem<20> ), .Y(n346) );
  OAI21X1 U550 ( .A(n936), .B(n944), .C(n347), .Y(n614) );
  OAI21X1 U551 ( .A(n8), .B(n943), .C(\mem<19> ), .Y(n347) );
  OAI21X1 U552 ( .A(n935), .B(n944), .C(n348), .Y(n615) );
  OAI21X1 U553 ( .A(n6), .B(n943), .C(\mem<18> ), .Y(n348) );
  OAI21X1 U554 ( .A(n934), .B(n944), .C(n349), .Y(n616) );
  OAI21X1 U555 ( .A(n4), .B(n943), .C(\mem<17> ), .Y(n349) );
  OAI21X1 U556 ( .A(n928), .B(n944), .C(n350), .Y(n617) );
  OAI21X1 U557 ( .A(n2), .B(n943), .C(\mem<16> ), .Y(n350) );
  OAI21X1 U561 ( .A(n81), .B(n933), .C(n352), .Y(n618) );
  OAI21X1 U562 ( .A(n32), .B(n929), .C(\mem<15> ), .Y(n352) );
  OAI21X1 U565 ( .A(n78), .B(n933), .C(n357), .Y(n619) );
  OAI21X1 U566 ( .A(n30), .B(n929), .C(\mem<14> ), .Y(n357) );
  OAI21X1 U569 ( .A(n942), .B(n933), .C(n359), .Y(n620) );
  OAI21X1 U570 ( .A(n28), .B(n929), .C(\mem<13> ), .Y(n359) );
  OAI21X1 U573 ( .A(n941), .B(n933), .C(n361), .Y(n621) );
  OAI21X1 U574 ( .A(n26), .B(n929), .C(\mem<12> ), .Y(n361) );
  OAI21X1 U577 ( .A(n75), .B(n933), .C(n363), .Y(n622) );
  OAI21X1 U578 ( .A(n24), .B(n929), .C(\mem<11> ), .Y(n363) );
  OAI21X1 U581 ( .A(n72), .B(n933), .C(n365), .Y(n623) );
  OAI21X1 U582 ( .A(n22), .B(n929), .C(\mem<10> ), .Y(n365) );
  OAI21X1 U585 ( .A(n69), .B(n933), .C(n366), .Y(n624) );
  OAI21X1 U586 ( .A(n20), .B(n929), .C(\mem<9> ), .Y(n366) );
  OAI21X1 U589 ( .A(n66), .B(n933), .C(n367), .Y(n625) );
  OAI21X1 U590 ( .A(n18), .B(n929), .C(\mem<8> ), .Y(n367) );
  OAI21X1 U593 ( .A(n940), .B(n932), .C(n368), .Y(n626) );
  OAI21X1 U594 ( .A(n16), .B(n929), .C(\mem<7> ), .Y(n368) );
  OAI21X1 U597 ( .A(n939), .B(n932), .C(n370), .Y(n627) );
  OAI21X1 U598 ( .A(n14), .B(n929), .C(\mem<6> ), .Y(n370) );
  OAI21X1 U601 ( .A(n938), .B(n932), .C(n371), .Y(n628) );
  OAI21X1 U602 ( .A(n12), .B(n929), .C(\mem<5> ), .Y(n371) );
  OAI21X1 U605 ( .A(n937), .B(n932), .C(n372), .Y(n629) );
  OAI21X1 U606 ( .A(n10), .B(n929), .C(\mem<4> ), .Y(n372) );
  OAI21X1 U610 ( .A(n936), .B(n932), .C(n373), .Y(n630) );
  OAI21X1 U611 ( .A(n8), .B(n929), .C(\mem<3> ), .Y(n373) );
  OAI21X1 U614 ( .A(n935), .B(n932), .C(n375), .Y(n631) );
  OAI21X1 U615 ( .A(n6), .B(n929), .C(\mem<2> ), .Y(n375) );
  OAI21X1 U618 ( .A(n934), .B(n932), .C(n376), .Y(n632) );
  OAI21X1 U619 ( .A(n4), .B(n929), .C(\mem<1> ), .Y(n376) );
  OAI21X1 U623 ( .A(n928), .B(n932), .C(n377), .Y(n633) );
  OAI21X1 U624 ( .A(n2), .B(n929), .C(\mem<0> ), .Y(n377) );
  NOR3X1 U634 ( .A(rst), .B(write), .C(n1003), .Y(data_out) );
  INVX4 U2 ( .A(n997), .Y(n996) );
  INVX8 U3 ( .A(n996), .Y(n916) );
  INVX2 U4 ( .A(n996), .Y(n915) );
  OR2X2 U5 ( .A(n997), .B(n998), .Y(n636) );
  AND2X2 U8 ( .A(n998), .B(n997), .Y(n358) );
  INVX1 U9 ( .A(N28), .Y(n1003) );
  INVX2 U10 ( .A(n916), .Y(n920) );
  INVX2 U11 ( .A(n916), .Y(n922) );
  INVX2 U12 ( .A(n916), .Y(n917) );
  INVX2 U13 ( .A(n908), .Y(n914) );
  INVX2 U14 ( .A(n908), .Y(n910) );
  INVX2 U15 ( .A(n908), .Y(n909) );
  INVX2 U16 ( .A(n916), .Y(n921) );
  INVX1 U17 ( .A(n1000), .Y(n906) );
  INVX1 U18 ( .A(n1000), .Y(n907) );
  INVX1 U19 ( .A(n902), .Y(n903) );
  INVX1 U20 ( .A(n902), .Y(n904) );
  AND2X1 U21 ( .A(N25), .B(n1005), .Y(n168) );
  INVX1 U22 ( .A(N24), .Y(n1005) );
  INVX1 U23 ( .A(N22), .Y(n1002) );
  AND2X1 U24 ( .A(data_in), .B(n931), .Y(n90) );
  AND2X1 U25 ( .A(N25), .B(N24), .Y(n91) );
  BUFX2 U26 ( .A(n90), .Y(n995) );
  AND2X1 U27 ( .A(N23), .B(n1001), .Y(n92) );
  AND2X1 U28 ( .A(N23), .B(n1002), .Y(n111) );
  AND2X1 U29 ( .A(n998), .B(n996), .Y(n356) );
  BUFX2 U30 ( .A(n90), .Y(n994) );
  BUFX2 U31 ( .A(n60), .Y(n931) );
  BUFX2 U32 ( .A(n60), .Y(n930) );
  BUFX2 U33 ( .A(n362), .Y(n993) );
  BUFX2 U34 ( .A(n354), .Y(n990) );
  BUFX2 U35 ( .A(n362), .Y(n992) );
  BUFX2 U36 ( .A(n351), .Y(n989) );
  BUFX2 U37 ( .A(n317), .Y(n986) );
  BUFX2 U38 ( .A(n351), .Y(n988) );
  BUFX2 U39 ( .A(n315), .Y(n985) );
  BUFX2 U40 ( .A(n315), .Y(n984) );
  BUFX2 U41 ( .A(n298), .Y(n982) );
  BUFX2 U42 ( .A(n298), .Y(n981) );
  BUFX2 U43 ( .A(n280), .Y(n979) );
  BUFX2 U44 ( .A(n262), .Y(n976) );
  BUFX2 U45 ( .A(n280), .Y(n978) );
  BUFX2 U46 ( .A(n244), .Y(n975) );
  BUFX2 U47 ( .A(n241), .Y(n972) );
  BUFX2 U48 ( .A(n244), .Y(n974) );
  BUFX2 U81 ( .A(n223), .Y(n971) );
  BUFX2 U82 ( .A(n205), .Y(n968) );
  BUFX2 U115 ( .A(n223), .Y(n970) );
  BUFX2 U116 ( .A(n187), .Y(n967) );
  BUFX2 U149 ( .A(n169), .Y(n964) );
  BUFX2 U150 ( .A(n187), .Y(n966) );
  BUFX2 U183 ( .A(n150), .Y(n963) );
  BUFX2 U184 ( .A(n150), .Y(n962) );
  BUFX2 U217 ( .A(n133), .Y(n960) );
  BUFX2 U218 ( .A(n133), .Y(n959) );
  BUFX2 U251 ( .A(n130), .Y(n957) );
  BUFX2 U252 ( .A(n130), .Y(n956) );
  BUFX2 U285 ( .A(n112), .Y(n954) );
  BUFX2 U286 ( .A(n112), .Y(n953) );
  BUFX2 U319 ( .A(n93), .Y(n951) );
  BUFX2 U320 ( .A(n93), .Y(n950) );
  BUFX2 U353 ( .A(n87), .Y(n948) );
  BUFX2 U354 ( .A(n87), .Y(n947) );
  BUFX2 U387 ( .A(n84), .Y(n945) );
  BUFX2 U388 ( .A(n84), .Y(n944) );
  BUFX2 U421 ( .A(n63), .Y(n933) );
  BUFX2 U422 ( .A(n63), .Y(n932) );
  INVX1 U455 ( .A(n999), .Y(n998) );
  INVX1 U456 ( .A(n998), .Y(n908) );
  INVX1 U457 ( .A(n34), .Y(n929) );
  INVX1 U490 ( .A(n45), .Y(n943) );
  INVX1 U491 ( .A(n50), .Y(n952) );
  INVX1 U524 ( .A(n51), .Y(n955) );
  INVX1 U525 ( .A(n56), .Y(n980) );
  INVX1 U558 ( .A(n57), .Y(n983) );
  INVX1 U559 ( .A(n1000), .Y(n905) );
  INVX1 U560 ( .A(n47), .Y(n946) );
  INVX1 U563 ( .A(n53), .Y(n958) );
  INVX1 U564 ( .A(n43), .Y(n941) );
  INVX1 U567 ( .A(n44), .Y(n942) );
  INVX1 U568 ( .A(n36), .Y(n935) );
  INVX1 U571 ( .A(n40), .Y(n939) );
  INVX1 U572 ( .A(n48), .Y(n949) );
  INVX1 U575 ( .A(n54), .Y(n961) );
  BUFX2 U576 ( .A(n169), .Y(n965) );
  BUFX2 U579 ( .A(n205), .Y(n969) );
  BUFX2 U580 ( .A(n241), .Y(n973) );
  BUFX2 U583 ( .A(n262), .Y(n977) );
  BUFX2 U584 ( .A(n317), .Y(n987) );
  BUFX2 U587 ( .A(n354), .Y(n991) );
  INVX1 U588 ( .A(n33), .Y(n928) );
  INVX1 U591 ( .A(n35), .Y(n934) );
  INVX1 U592 ( .A(n37), .Y(n936) );
  INVX1 U595 ( .A(n38), .Y(n937) );
  INVX1 U596 ( .A(n39), .Y(n938) );
  INVX1 U599 ( .A(n41), .Y(n940) );
  INVX1 U600 ( .A(n1002), .Y(n1001) );
  OR2X2 U603 ( .A(n1000), .B(N21), .Y(n644) );
  OR2X2 U604 ( .A(n905), .B(N21), .Y(n640) );
  INVX1 U607 ( .A(N21), .Y(n902) );
  INVX1 U608 ( .A(write), .Y(n1004) );
  AND2X1 U609 ( .A(n33), .B(n930), .Y(n1) );
  INVX1 U612 ( .A(n1), .Y(n2) );
  AND2X1 U613 ( .A(n35), .B(n930), .Y(n3) );
  INVX1 U616 ( .A(n3), .Y(n4) );
  AND2X1 U617 ( .A(n36), .B(n930), .Y(n5) );
  INVX1 U620 ( .A(n5), .Y(n6) );
  AND2X1 U621 ( .A(n37), .B(n930), .Y(n7) );
  INVX1 U622 ( .A(n7), .Y(n8) );
  AND2X1 U625 ( .A(n38), .B(n930), .Y(n9) );
  INVX1 U626 ( .A(n9), .Y(n10) );
  AND2X1 U627 ( .A(n39), .B(n930), .Y(n11) );
  INVX1 U628 ( .A(n11), .Y(n12) );
  AND2X1 U629 ( .A(n40), .B(n930), .Y(n13) );
  INVX1 U630 ( .A(n13), .Y(n14) );
  AND2X1 U631 ( .A(n41), .B(n930), .Y(n15) );
  INVX1 U632 ( .A(n15), .Y(n16) );
  AND2X1 U633 ( .A(n65), .B(n931), .Y(n17) );
  INVX1 U635 ( .A(n17), .Y(n18) );
  AND2X1 U636 ( .A(n68), .B(n931), .Y(n19) );
  INVX1 U637 ( .A(n19), .Y(n20) );
  AND2X1 U638 ( .A(n71), .B(n931), .Y(n21) );
  INVX1 U639 ( .A(n21), .Y(n22) );
  AND2X1 U640 ( .A(n74), .B(n931), .Y(n23) );
  INVX1 U641 ( .A(n23), .Y(n24) );
  AND2X1 U642 ( .A(n43), .B(n931), .Y(n25) );
  INVX1 U643 ( .A(n25), .Y(n26) );
  AND2X1 U644 ( .A(n44), .B(n931), .Y(n27) );
  INVX1 U645 ( .A(n27), .Y(n28) );
  AND2X1 U646 ( .A(n77), .B(n931), .Y(n29) );
  INVX1 U647 ( .A(n29), .Y(n30) );
  AND2X1 U648 ( .A(n80), .B(n931), .Y(n31) );
  INVX1 U649 ( .A(n31), .Y(n32) );
  AND2X1 U650 ( .A(n641), .B(n374), .Y(n33) );
  AND2X1 U651 ( .A(n643), .B(n635), .Y(n34) );
  AND2X1 U652 ( .A(n641), .B(n637), .Y(n35) );
  AND2X1 U653 ( .A(n641), .B(n358), .Y(n36) );
  AND2X1 U654 ( .A(n641), .B(n356), .Y(n37) );
  AND2X1 U655 ( .A(n645), .B(n374), .Y(n38) );
  AND2X1 U656 ( .A(n645), .B(n637), .Y(n39) );
  AND2X1 U657 ( .A(n645), .B(n358), .Y(n40) );
  AND2X1 U658 ( .A(n645), .B(n356), .Y(n41) );
  AND2X1 U659 ( .A(n374), .B(n355), .Y(n43) );
  AND2X1 U660 ( .A(n637), .B(n355), .Y(n44) );
  AND2X1 U661 ( .A(n643), .B(n639), .Y(n45) );
  AND2X1 U662 ( .A(n643), .B(n111), .Y(n47) );
  AND2X1 U663 ( .A(n643), .B(n92), .Y(n48) );
  AND2X1 U664 ( .A(n647), .B(n635), .Y(n50) );
  AND2X1 U665 ( .A(n647), .B(n639), .Y(n51) );
  AND2X1 U666 ( .A(n647), .B(n111), .Y(n53) );
  AND2X1 U667 ( .A(n647), .B(n92), .Y(n54) );
  AND2X1 U668 ( .A(n635), .B(n91), .Y(n56) );
  AND2X1 U669 ( .A(n639), .B(n91), .Y(n57) );
  OR2X1 U670 ( .A(n1004), .B(rst), .Y(n59) );
  INVX1 U671 ( .A(n59), .Y(n60) );
  AND2X1 U672 ( .A(n34), .B(n994), .Y(n62) );
  INVX1 U673 ( .A(n62), .Y(n63) );
  AND2X1 U674 ( .A(n364), .B(n374), .Y(n65) );
  INVX1 U675 ( .A(n65), .Y(n66) );
  AND2X1 U676 ( .A(n364), .B(n637), .Y(n68) );
  INVX1 U677 ( .A(n68), .Y(n69) );
  AND2X1 U678 ( .A(n364), .B(n358), .Y(n71) );
  INVX1 U679 ( .A(n71), .Y(n72) );
  AND2X1 U680 ( .A(n364), .B(n356), .Y(n74) );
  INVX1 U681 ( .A(n74), .Y(n75) );
  AND2X1 U682 ( .A(n358), .B(n355), .Y(n77) );
  INVX1 U683 ( .A(n77), .Y(n78) );
  AND2X1 U684 ( .A(n355), .B(n356), .Y(n80) );
  INVX1 U685 ( .A(n80), .Y(n81) );
  AND2X1 U686 ( .A(n45), .B(n994), .Y(n83) );
  INVX1 U687 ( .A(n83), .Y(n84) );
  AND2X1 U688 ( .A(n47), .B(n994), .Y(n86) );
  INVX1 U689 ( .A(n86), .Y(n87) );
  AND2X1 U690 ( .A(n48), .B(n994), .Y(n89) );
  INVX1 U691 ( .A(n89), .Y(n93) );
  AND2X1 U692 ( .A(n50), .B(n994), .Y(n95) );
  INVX1 U693 ( .A(n95), .Y(n112) );
  AND2X1 U694 ( .A(n51), .B(n994), .Y(n114) );
  INVX1 U695 ( .A(n114), .Y(n130) );
  AND2X1 U696 ( .A(n53), .B(n994), .Y(n131) );
  INVX1 U697 ( .A(n131), .Y(n133) );
  AND2X1 U698 ( .A(n54), .B(n995), .Y(n149) );
  INVX1 U699 ( .A(n149), .Y(n150) );
  AND2X1 U700 ( .A(n168), .B(n635), .Y(n152) );
  INVX1 U701 ( .A(n152), .Y(n169) );
  AND2X1 U702 ( .A(n152), .B(n995), .Y(n171) );
  INVX1 U703 ( .A(n171), .Y(n187) );
  AND2X1 U704 ( .A(n168), .B(n639), .Y(n189) );
  INVX1 U705 ( .A(n189), .Y(n205) );
  AND2X1 U706 ( .A(n189), .B(n995), .Y(n207) );
  INVX1 U707 ( .A(n207), .Y(n223) );
  AND2X1 U708 ( .A(n168), .B(n111), .Y(n225) );
  INVX1 U709 ( .A(n225), .Y(n241) );
  AND2X1 U710 ( .A(n225), .B(n995), .Y(n242) );
  INVX1 U711 ( .A(n242), .Y(n244) );
  AND2X1 U712 ( .A(n168), .B(n92), .Y(n260) );
  INVX1 U713 ( .A(n260), .Y(n262) );
  AND2X1 U714 ( .A(n260), .B(n995), .Y(n278) );
  INVX1 U715 ( .A(n278), .Y(n280) );
  AND2X1 U716 ( .A(n56), .B(n995), .Y(n296) );
  INVX1 U717 ( .A(n296), .Y(n298) );
  AND2X1 U718 ( .A(n57), .B(n995), .Y(n314) );
  INVX1 U719 ( .A(n314), .Y(n315) );
  INVX1 U720 ( .A(n333), .Y(n317) );
  AND2X1 U721 ( .A(n111), .B(n91), .Y(n333) );
  AND2X1 U722 ( .A(n333), .B(n995), .Y(n335) );
  INVX1 U723 ( .A(n335), .Y(n351) );
  AND2X1 U724 ( .A(n91), .B(n92), .Y(n353) );
  INVX1 U725 ( .A(n353), .Y(n354) );
  AND2X1 U726 ( .A(n994), .B(n353), .Y(n360) );
  INVX1 U727 ( .A(n360), .Y(n362) );
  OR2X1 U728 ( .A(n996), .B(n998), .Y(n369) );
  INVX1 U729 ( .A(n369), .Y(n374) );
  OR2X1 U730 ( .A(n1001), .B(N23), .Y(n634) );
  INVX1 U731 ( .A(n634), .Y(n635) );
  INVX1 U732 ( .A(n636), .Y(n637) );
  OR2X1 U733 ( .A(n1002), .B(N23), .Y(n638) );
  INVX1 U734 ( .A(n638), .Y(n639) );
  INVX1 U735 ( .A(n640), .Y(n641) );
  OR2X1 U736 ( .A(N24), .B(N25), .Y(n642) );
  INVX1 U737 ( .A(n642), .Y(n643) );
  INVX1 U738 ( .A(n644), .Y(n645) );
  OR2X1 U739 ( .A(n1005), .B(N25), .Y(n646) );
  INVX1 U740 ( .A(n646), .Y(n647) );
  MUX2X1 U741 ( .B(n649), .A(n650), .S(n914), .Y(n648) );
  MUX2X1 U742 ( .B(n652), .A(n653), .S(n914), .Y(n651) );
  MUX2X1 U743 ( .B(n655), .A(n656), .S(n914), .Y(n654) );
  MUX2X1 U744 ( .B(n658), .A(n659), .S(n914), .Y(n657) );
  MUX2X1 U745 ( .B(n661), .A(n662), .S(n904), .Y(n660) );
  MUX2X1 U746 ( .B(n664), .A(n665), .S(n914), .Y(n663) );
  MUX2X1 U747 ( .B(n667), .A(n668), .S(n914), .Y(n666) );
  MUX2X1 U748 ( .B(n670), .A(n671), .S(n914), .Y(n669) );
  MUX2X1 U749 ( .B(n673), .A(n674), .S(n914), .Y(n672) );
  MUX2X1 U750 ( .B(n676), .A(n677), .S(n904), .Y(n675) );
  MUX2X1 U751 ( .B(n679), .A(n680), .S(n914), .Y(n678) );
  MUX2X1 U752 ( .B(n682), .A(n683), .S(n914), .Y(n681) );
  MUX2X1 U753 ( .B(n685), .A(n686), .S(n914), .Y(n684) );
  MUX2X1 U754 ( .B(n688), .A(n689), .S(n914), .Y(n687) );
  MUX2X1 U755 ( .B(n691), .A(n692), .S(n904), .Y(n690) );
  MUX2X1 U756 ( .B(n694), .A(n695), .S(n913), .Y(n693) );
  MUX2X1 U757 ( .B(n697), .A(n698), .S(n913), .Y(n696) );
  MUX2X1 U758 ( .B(n700), .A(n701), .S(n913), .Y(n699) );
  MUX2X1 U759 ( .B(n703), .A(n704), .S(n913), .Y(n702) );
  MUX2X1 U760 ( .B(n706), .A(n707), .S(n904), .Y(n705) );
  MUX2X1 U761 ( .B(n709), .A(n710), .S(N23), .Y(n708) );
  MUX2X1 U762 ( .B(n712), .A(n713), .S(n913), .Y(n711) );
  MUX2X1 U763 ( .B(n715), .A(n716), .S(n913), .Y(n714) );
  MUX2X1 U764 ( .B(n718), .A(n719), .S(n913), .Y(n717) );
  MUX2X1 U765 ( .B(n721), .A(n722), .S(n913), .Y(n720) );
  MUX2X1 U766 ( .B(n724), .A(n725), .S(n904), .Y(n723) );
  MUX2X1 U767 ( .B(n727), .A(n728), .S(n913), .Y(n726) );
  MUX2X1 U768 ( .B(n730), .A(n731), .S(n913), .Y(n729) );
  MUX2X1 U769 ( .B(n733), .A(n734), .S(n913), .Y(n732) );
  MUX2X1 U770 ( .B(n736), .A(n737), .S(n913), .Y(n735) );
  MUX2X1 U771 ( .B(n739), .A(n740), .S(n904), .Y(n738) );
  MUX2X1 U772 ( .B(n742), .A(n743), .S(n912), .Y(n741) );
  MUX2X1 U773 ( .B(n745), .A(n746), .S(n912), .Y(n744) );
  MUX2X1 U774 ( .B(n748), .A(n749), .S(n912), .Y(n747) );
  MUX2X1 U775 ( .B(n751), .A(n752), .S(n912), .Y(n750) );
  MUX2X1 U776 ( .B(n754), .A(n755), .S(n904), .Y(n753) );
  MUX2X1 U777 ( .B(n757), .A(n758), .S(n912), .Y(n756) );
  MUX2X1 U778 ( .B(n760), .A(n761), .S(n912), .Y(n759) );
  MUX2X1 U779 ( .B(n763), .A(n764), .S(n912), .Y(n762) );
  MUX2X1 U780 ( .B(n766), .A(n767), .S(n912), .Y(n765) );
  MUX2X1 U781 ( .B(n769), .A(n770), .S(n904), .Y(n768) );
  MUX2X1 U782 ( .B(n772), .A(n773), .S(N23), .Y(n771) );
  MUX2X1 U783 ( .B(n775), .A(n776), .S(n912), .Y(n774) );
  MUX2X1 U784 ( .B(n778), .A(n779), .S(n912), .Y(n777) );
  MUX2X1 U785 ( .B(n781), .A(n782), .S(n912), .Y(n780) );
  MUX2X1 U786 ( .B(n784), .A(n785), .S(n912), .Y(n783) );
  MUX2X1 U787 ( .B(n787), .A(n788), .S(n904), .Y(n786) );
  MUX2X1 U788 ( .B(n790), .A(n791), .S(n911), .Y(n789) );
  MUX2X1 U789 ( .B(n793), .A(n794), .S(n911), .Y(n792) );
  MUX2X1 U790 ( .B(n796), .A(n797), .S(n911), .Y(n795) );
  MUX2X1 U791 ( .B(n799), .A(n800), .S(n911), .Y(n798) );
  MUX2X1 U792 ( .B(n802), .A(n803), .S(n904), .Y(n801) );
  MUX2X1 U793 ( .B(n805), .A(n806), .S(n911), .Y(n804) );
  MUX2X1 U794 ( .B(n808), .A(n809), .S(n911), .Y(n807) );
  MUX2X1 U795 ( .B(n811), .A(n812), .S(n911), .Y(n810) );
  MUX2X1 U796 ( .B(n814), .A(n815), .S(n911), .Y(n813) );
  MUX2X1 U797 ( .B(n817), .A(n818), .S(n904), .Y(n816) );
  MUX2X1 U798 ( .B(n820), .A(n821), .S(n911), .Y(n819) );
  MUX2X1 U799 ( .B(n823), .A(n824), .S(n911), .Y(n822) );
  MUX2X1 U800 ( .B(n826), .A(n827), .S(n911), .Y(n825) );
  MUX2X1 U801 ( .B(n829), .A(n830), .S(n911), .Y(n828) );
  MUX2X1 U802 ( .B(n832), .A(n833), .S(n904), .Y(n831) );
  MUX2X1 U803 ( .B(n835), .A(n836), .S(N23), .Y(n834) );
  MUX2X1 U804 ( .B(n838), .A(n839), .S(n910), .Y(n837) );
  MUX2X1 U805 ( .B(n841), .A(n842), .S(n910), .Y(n840) );
  MUX2X1 U806 ( .B(n844), .A(n845), .S(n910), .Y(n843) );
  MUX2X1 U807 ( .B(n847), .A(n848), .S(n910), .Y(n846) );
  MUX2X1 U808 ( .B(n850), .A(n851), .S(n903), .Y(n849) );
  MUX2X1 U809 ( .B(n853), .A(n854), .S(n910), .Y(n852) );
  MUX2X1 U810 ( .B(n856), .A(n857), .S(n910), .Y(n855) );
  MUX2X1 U811 ( .B(n859), .A(n860), .S(n910), .Y(n858) );
  MUX2X1 U812 ( .B(n862), .A(n863), .S(n910), .Y(n861) );
  MUX2X1 U813 ( .B(n865), .A(n866), .S(n903), .Y(n864) );
  MUX2X1 U814 ( .B(n868), .A(n869), .S(n910), .Y(n867) );
  MUX2X1 U815 ( .B(n871), .A(n872), .S(n910), .Y(n870) );
  MUX2X1 U816 ( .B(n874), .A(n875), .S(n910), .Y(n873) );
  MUX2X1 U817 ( .B(n877), .A(n878), .S(n910), .Y(n876) );
  MUX2X1 U818 ( .B(n880), .A(n881), .S(n903), .Y(n879) );
  MUX2X1 U819 ( .B(n883), .A(n884), .S(n909), .Y(n882) );
  MUX2X1 U820 ( .B(n886), .A(n887), .S(n909), .Y(n885) );
  MUX2X1 U821 ( .B(n889), .A(n890), .S(n909), .Y(n888) );
  MUX2X1 U822 ( .B(n892), .A(n893), .S(n909), .Y(n891) );
  MUX2X1 U823 ( .B(n895), .A(n896), .S(n903), .Y(n894) );
  MUX2X1 U824 ( .B(n898), .A(n899), .S(N23), .Y(n897) );
  MUX2X1 U825 ( .B(n900), .A(n901), .S(N25), .Y(N28) );
  MUX2X1 U826 ( .B(\mem<254> ), .A(\mem<255> ), .S(n917), .Y(n650) );
  MUX2X1 U827 ( .B(\mem<252> ), .A(\mem<253> ), .S(n917), .Y(n649) );
  MUX2X1 U828 ( .B(\mem<250> ), .A(\mem<251> ), .S(n917), .Y(n653) );
  MUX2X1 U829 ( .B(\mem<248> ), .A(\mem<249> ), .S(n917), .Y(n652) );
  MUX2X1 U830 ( .B(n651), .A(n648), .S(n907), .Y(n662) );
  MUX2X1 U831 ( .B(\mem<246> ), .A(\mem<247> ), .S(n917), .Y(n656) );
  MUX2X1 U832 ( .B(\mem<244> ), .A(\mem<245> ), .S(n917), .Y(n655) );
  MUX2X1 U833 ( .B(\mem<242> ), .A(\mem<243> ), .S(n917), .Y(n659) );
  MUX2X1 U834 ( .B(\mem<240> ), .A(\mem<241> ), .S(n917), .Y(n658) );
  MUX2X1 U835 ( .B(n657), .A(n654), .S(n907), .Y(n661) );
  MUX2X1 U836 ( .B(\mem<238> ), .A(\mem<239> ), .S(n918), .Y(n665) );
  MUX2X1 U837 ( .B(\mem<236> ), .A(\mem<237> ), .S(n918), .Y(n664) );
  MUX2X1 U838 ( .B(\mem<234> ), .A(\mem<235> ), .S(n918), .Y(n668) );
  MUX2X1 U839 ( .B(\mem<232> ), .A(\mem<233> ), .S(n918), .Y(n667) );
  MUX2X1 U840 ( .B(n666), .A(n663), .S(n907), .Y(n677) );
  MUX2X1 U841 ( .B(\mem<230> ), .A(\mem<231> ), .S(n918), .Y(n671) );
  MUX2X1 U842 ( .B(\mem<228> ), .A(\mem<229> ), .S(n918), .Y(n670) );
  MUX2X1 U843 ( .B(\mem<226> ), .A(\mem<227> ), .S(n918), .Y(n674) );
  MUX2X1 U844 ( .B(\mem<224> ), .A(\mem<225> ), .S(n918), .Y(n673) );
  MUX2X1 U845 ( .B(n672), .A(n669), .S(n907), .Y(n676) );
  MUX2X1 U846 ( .B(n675), .A(n660), .S(n1001), .Y(n710) );
  MUX2X1 U847 ( .B(\mem<222> ), .A(\mem<223> ), .S(n918), .Y(n680) );
  MUX2X1 U848 ( .B(\mem<220> ), .A(\mem<221> ), .S(n918), .Y(n679) );
  MUX2X1 U849 ( .B(\mem<218> ), .A(\mem<219> ), .S(n918), .Y(n683) );
  MUX2X1 U850 ( .B(\mem<216> ), .A(\mem<217> ), .S(n918), .Y(n682) );
  MUX2X1 U851 ( .B(n681), .A(n678), .S(n907), .Y(n692) );
  MUX2X1 U852 ( .B(\mem<214> ), .A(\mem<215> ), .S(n919), .Y(n686) );
  MUX2X1 U853 ( .B(\mem<212> ), .A(\mem<213> ), .S(n919), .Y(n685) );
  MUX2X1 U854 ( .B(\mem<210> ), .A(\mem<211> ), .S(n919), .Y(n689) );
  MUX2X1 U855 ( .B(\mem<208> ), .A(\mem<209> ), .S(n919), .Y(n688) );
  MUX2X1 U856 ( .B(n687), .A(n684), .S(n907), .Y(n691) );
  MUX2X1 U857 ( .B(\mem<206> ), .A(\mem<207> ), .S(n919), .Y(n695) );
  MUX2X1 U858 ( .B(\mem<204> ), .A(\mem<205> ), .S(n919), .Y(n694) );
  MUX2X1 U859 ( .B(\mem<202> ), .A(\mem<203> ), .S(n919), .Y(n698) );
  MUX2X1 U860 ( .B(\mem<200> ), .A(\mem<201> ), .S(n919), .Y(n697) );
  MUX2X1 U861 ( .B(n696), .A(n693), .S(n907), .Y(n707) );
  MUX2X1 U862 ( .B(\mem<198> ), .A(\mem<199> ), .S(n919), .Y(n701) );
  MUX2X1 U863 ( .B(\mem<196> ), .A(\mem<197> ), .S(n919), .Y(n700) );
  MUX2X1 U864 ( .B(\mem<194> ), .A(\mem<195> ), .S(n919), .Y(n704) );
  MUX2X1 U865 ( .B(\mem<192> ), .A(\mem<193> ), .S(n919), .Y(n703) );
  MUX2X1 U866 ( .B(n702), .A(n699), .S(n907), .Y(n706) );
  MUX2X1 U867 ( .B(n705), .A(n690), .S(n1001), .Y(n709) );
  MUX2X1 U868 ( .B(\mem<190> ), .A(\mem<191> ), .S(n920), .Y(n713) );
  MUX2X1 U869 ( .B(\mem<188> ), .A(\mem<189> ), .S(n920), .Y(n712) );
  MUX2X1 U870 ( .B(\mem<186> ), .A(\mem<187> ), .S(n920), .Y(n716) );
  MUX2X1 U871 ( .B(\mem<184> ), .A(\mem<185> ), .S(n920), .Y(n715) );
  MUX2X1 U872 ( .B(n714), .A(n711), .S(n907), .Y(n725) );
  MUX2X1 U873 ( .B(\mem<182> ), .A(\mem<183> ), .S(n920), .Y(n719) );
  MUX2X1 U874 ( .B(\mem<180> ), .A(\mem<181> ), .S(n920), .Y(n718) );
  MUX2X1 U875 ( .B(\mem<178> ), .A(\mem<179> ), .S(n920), .Y(n722) );
  MUX2X1 U876 ( .B(\mem<176> ), .A(\mem<177> ), .S(n920), .Y(n721) );
  MUX2X1 U877 ( .B(n720), .A(n717), .S(n907), .Y(n724) );
  MUX2X1 U878 ( .B(\mem<174> ), .A(\mem<175> ), .S(n920), .Y(n728) );
  MUX2X1 U879 ( .B(\mem<172> ), .A(\mem<173> ), .S(n920), .Y(n727) );
  MUX2X1 U880 ( .B(\mem<170> ), .A(\mem<171> ), .S(n920), .Y(n731) );
  MUX2X1 U881 ( .B(\mem<168> ), .A(\mem<169> ), .S(n920), .Y(n730) );
  MUX2X1 U882 ( .B(n729), .A(n726), .S(n907), .Y(n740) );
  MUX2X1 U883 ( .B(\mem<166> ), .A(\mem<167> ), .S(n921), .Y(n734) );
  MUX2X1 U884 ( .B(\mem<164> ), .A(\mem<165> ), .S(n921), .Y(n733) );
  MUX2X1 U885 ( .B(\mem<162> ), .A(\mem<163> ), .S(n921), .Y(n737) );
  MUX2X1 U886 ( .B(\mem<160> ), .A(\mem<161> ), .S(n921), .Y(n736) );
  MUX2X1 U887 ( .B(n735), .A(n732), .S(n907), .Y(n739) );
  MUX2X1 U888 ( .B(n738), .A(n723), .S(n1001), .Y(n773) );
  MUX2X1 U889 ( .B(\mem<158> ), .A(\mem<159> ), .S(n921), .Y(n743) );
  MUX2X1 U890 ( .B(\mem<156> ), .A(\mem<157> ), .S(n921), .Y(n742) );
  MUX2X1 U891 ( .B(\mem<154> ), .A(\mem<155> ), .S(n921), .Y(n746) );
  MUX2X1 U892 ( .B(\mem<152> ), .A(\mem<153> ), .S(n921), .Y(n745) );
  MUX2X1 U893 ( .B(n744), .A(n741), .S(n906), .Y(n755) );
  MUX2X1 U894 ( .B(\mem<150> ), .A(\mem<151> ), .S(n921), .Y(n749) );
  MUX2X1 U895 ( .B(\mem<148> ), .A(\mem<149> ), .S(n921), .Y(n748) );
  MUX2X1 U896 ( .B(\mem<146> ), .A(\mem<147> ), .S(n921), .Y(n752) );
  MUX2X1 U897 ( .B(\mem<144> ), .A(\mem<145> ), .S(n921), .Y(n751) );
  MUX2X1 U898 ( .B(n750), .A(n747), .S(n906), .Y(n754) );
  MUX2X1 U899 ( .B(\mem<142> ), .A(\mem<143> ), .S(n922), .Y(n758) );
  MUX2X1 U900 ( .B(\mem<140> ), .A(\mem<141> ), .S(n922), .Y(n757) );
  MUX2X1 U901 ( .B(\mem<138> ), .A(\mem<139> ), .S(n922), .Y(n761) );
  MUX2X1 U902 ( .B(\mem<136> ), .A(\mem<137> ), .S(n922), .Y(n760) );
  MUX2X1 U903 ( .B(n759), .A(n756), .S(n906), .Y(n770) );
  MUX2X1 U904 ( .B(\mem<134> ), .A(\mem<135> ), .S(n922), .Y(n764) );
  MUX2X1 U905 ( .B(\mem<132> ), .A(\mem<133> ), .S(n922), .Y(n763) );
  MUX2X1 U906 ( .B(\mem<130> ), .A(\mem<131> ), .S(n922), .Y(n767) );
  MUX2X1 U907 ( .B(\mem<128> ), .A(\mem<129> ), .S(n922), .Y(n766) );
  MUX2X1 U908 ( .B(n765), .A(n762), .S(n906), .Y(n769) );
  MUX2X1 U909 ( .B(n768), .A(n753), .S(n1001), .Y(n772) );
  MUX2X1 U910 ( .B(n771), .A(n708), .S(N24), .Y(n901) );
  MUX2X1 U911 ( .B(\mem<126> ), .A(\mem<127> ), .S(n922), .Y(n776) );
  MUX2X1 U912 ( .B(\mem<124> ), .A(\mem<125> ), .S(n922), .Y(n775) );
  MUX2X1 U913 ( .B(\mem<122> ), .A(\mem<123> ), .S(n922), .Y(n779) );
  MUX2X1 U914 ( .B(\mem<120> ), .A(\mem<121> ), .S(n922), .Y(n778) );
  MUX2X1 U915 ( .B(n777), .A(n774), .S(n906), .Y(n788) );
  MUX2X1 U916 ( .B(\mem<118> ), .A(\mem<119> ), .S(n923), .Y(n782) );
  MUX2X1 U917 ( .B(\mem<116> ), .A(\mem<117> ), .S(n923), .Y(n781) );
  MUX2X1 U918 ( .B(\mem<114> ), .A(\mem<115> ), .S(n923), .Y(n785) );
  MUX2X1 U919 ( .B(\mem<112> ), .A(\mem<113> ), .S(n923), .Y(n784) );
  MUX2X1 U920 ( .B(n783), .A(n780), .S(n906), .Y(n787) );
  MUX2X1 U921 ( .B(\mem<110> ), .A(\mem<111> ), .S(n923), .Y(n791) );
  MUX2X1 U922 ( .B(\mem<108> ), .A(\mem<109> ), .S(n923), .Y(n790) );
  MUX2X1 U923 ( .B(\mem<106> ), .A(\mem<107> ), .S(n923), .Y(n794) );
  MUX2X1 U924 ( .B(\mem<104> ), .A(\mem<105> ), .S(n923), .Y(n793) );
  MUX2X1 U925 ( .B(n792), .A(n789), .S(n906), .Y(n803) );
  MUX2X1 U926 ( .B(\mem<102> ), .A(\mem<103> ), .S(n923), .Y(n797) );
  MUX2X1 U927 ( .B(\mem<100> ), .A(\mem<101> ), .S(n923), .Y(n796) );
  MUX2X1 U928 ( .B(\mem<98> ), .A(\mem<99> ), .S(n923), .Y(n800) );
  MUX2X1 U929 ( .B(\mem<96> ), .A(\mem<97> ), .S(n923), .Y(n799) );
  MUX2X1 U930 ( .B(n798), .A(n795), .S(n906), .Y(n802) );
  MUX2X1 U931 ( .B(n801), .A(n786), .S(n1001), .Y(n836) );
  MUX2X1 U932 ( .B(\mem<94> ), .A(\mem<95> ), .S(n924), .Y(n806) );
  MUX2X1 U933 ( .B(\mem<92> ), .A(\mem<93> ), .S(n924), .Y(n805) );
  MUX2X1 U934 ( .B(\mem<90> ), .A(\mem<91> ), .S(n924), .Y(n809) );
  MUX2X1 U935 ( .B(\mem<88> ), .A(\mem<89> ), .S(n924), .Y(n808) );
  MUX2X1 U936 ( .B(n807), .A(n804), .S(n906), .Y(n818) );
  MUX2X1 U937 ( .B(\mem<86> ), .A(\mem<87> ), .S(n924), .Y(n812) );
  MUX2X1 U938 ( .B(\mem<84> ), .A(\mem<85> ), .S(n924), .Y(n811) );
  MUX2X1 U939 ( .B(\mem<82> ), .A(\mem<83> ), .S(n924), .Y(n815) );
  MUX2X1 U940 ( .B(\mem<80> ), .A(\mem<81> ), .S(n924), .Y(n814) );
  MUX2X1 U941 ( .B(n813), .A(n810), .S(n906), .Y(n817) );
  MUX2X1 U942 ( .B(\mem<78> ), .A(\mem<79> ), .S(n924), .Y(n821) );
  MUX2X1 U943 ( .B(\mem<76> ), .A(\mem<77> ), .S(n924), .Y(n820) );
  MUX2X1 U944 ( .B(\mem<74> ), .A(\mem<75> ), .S(n924), .Y(n824) );
  MUX2X1 U945 ( .B(\mem<72> ), .A(\mem<73> ), .S(n924), .Y(n823) );
  MUX2X1 U946 ( .B(n822), .A(n819), .S(n906), .Y(n833) );
  MUX2X1 U947 ( .B(\mem<70> ), .A(\mem<71> ), .S(n925), .Y(n827) );
  MUX2X1 U948 ( .B(\mem<68> ), .A(\mem<69> ), .S(n925), .Y(n826) );
  MUX2X1 U949 ( .B(\mem<66> ), .A(\mem<67> ), .S(n925), .Y(n830) );
  MUX2X1 U950 ( .B(\mem<64> ), .A(\mem<65> ), .S(n925), .Y(n829) );
  MUX2X1 U951 ( .B(n828), .A(n825), .S(n906), .Y(n832) );
  MUX2X1 U952 ( .B(n831), .A(n816), .S(n1001), .Y(n835) );
  MUX2X1 U953 ( .B(\mem<62> ), .A(\mem<63> ), .S(n925), .Y(n839) );
  MUX2X1 U954 ( .B(\mem<60> ), .A(\mem<61> ), .S(n925), .Y(n838) );
  MUX2X1 U955 ( .B(\mem<58> ), .A(\mem<59> ), .S(n925), .Y(n842) );
  MUX2X1 U956 ( .B(\mem<56> ), .A(\mem<57> ), .S(n925), .Y(n841) );
  MUX2X1 U957 ( .B(n840), .A(n837), .S(n905), .Y(n851) );
  MUX2X1 U958 ( .B(\mem<54> ), .A(\mem<55> ), .S(n925), .Y(n845) );
  MUX2X1 U959 ( .B(\mem<52> ), .A(\mem<53> ), .S(n925), .Y(n844) );
  MUX2X1 U960 ( .B(\mem<50> ), .A(\mem<51> ), .S(n925), .Y(n848) );
  MUX2X1 U961 ( .B(\mem<48> ), .A(\mem<49> ), .S(n925), .Y(n847) );
  MUX2X1 U962 ( .B(n846), .A(n843), .S(n905), .Y(n850) );
  MUX2X1 U963 ( .B(\mem<46> ), .A(\mem<47> ), .S(n926), .Y(n854) );
  MUX2X1 U964 ( .B(\mem<44> ), .A(\mem<45> ), .S(n926), .Y(n853) );
  MUX2X1 U965 ( .B(\mem<42> ), .A(\mem<43> ), .S(n926), .Y(n857) );
  MUX2X1 U966 ( .B(\mem<40> ), .A(\mem<41> ), .S(n926), .Y(n856) );
  MUX2X1 U967 ( .B(n855), .A(n852), .S(n905), .Y(n866) );
  MUX2X1 U968 ( .B(\mem<38> ), .A(\mem<39> ), .S(n926), .Y(n860) );
  MUX2X1 U969 ( .B(\mem<36> ), .A(\mem<37> ), .S(n926), .Y(n859) );
  MUX2X1 U970 ( .B(\mem<34> ), .A(\mem<35> ), .S(n926), .Y(n863) );
  MUX2X1 U971 ( .B(\mem<32> ), .A(\mem<33> ), .S(n926), .Y(n862) );
  MUX2X1 U972 ( .B(n861), .A(n858), .S(n905), .Y(n865) );
  MUX2X1 U973 ( .B(n864), .A(n849), .S(n1001), .Y(n899) );
  MUX2X1 U974 ( .B(\mem<30> ), .A(\mem<31> ), .S(n926), .Y(n869) );
  MUX2X1 U975 ( .B(\mem<28> ), .A(\mem<29> ), .S(n926), .Y(n868) );
  MUX2X1 U976 ( .B(\mem<26> ), .A(\mem<27> ), .S(n926), .Y(n872) );
  MUX2X1 U977 ( .B(\mem<24> ), .A(\mem<25> ), .S(n926), .Y(n871) );
  MUX2X1 U978 ( .B(n870), .A(n867), .S(n905), .Y(n881) );
  MUX2X1 U979 ( .B(\mem<22> ), .A(\mem<23> ), .S(n927), .Y(n875) );
  MUX2X1 U980 ( .B(\mem<20> ), .A(\mem<21> ), .S(n927), .Y(n874) );
  MUX2X1 U981 ( .B(\mem<18> ), .A(\mem<19> ), .S(n927), .Y(n878) );
  MUX2X1 U982 ( .B(\mem<16> ), .A(\mem<17> ), .S(n927), .Y(n877) );
  MUX2X1 U983 ( .B(n876), .A(n873), .S(n905), .Y(n880) );
  MUX2X1 U984 ( .B(\mem<14> ), .A(\mem<15> ), .S(n927), .Y(n884) );
  MUX2X1 U985 ( .B(\mem<12> ), .A(\mem<13> ), .S(n927), .Y(n883) );
  MUX2X1 U986 ( .B(\mem<10> ), .A(\mem<11> ), .S(n927), .Y(n887) );
  MUX2X1 U987 ( .B(\mem<8> ), .A(\mem<9> ), .S(n927), .Y(n886) );
  MUX2X1 U988 ( .B(n885), .A(n882), .S(n905), .Y(n896) );
  MUX2X1 U989 ( .B(\mem<6> ), .A(\mem<7> ), .S(n927), .Y(n890) );
  MUX2X1 U990 ( .B(\mem<4> ), .A(\mem<5> ), .S(n927), .Y(n889) );
  MUX2X1 U991 ( .B(\mem<2> ), .A(\mem<3> ), .S(n927), .Y(n893) );
  MUX2X1 U992 ( .B(\mem<0> ), .A(\mem<1> ), .S(n927), .Y(n892) );
  MUX2X1 U993 ( .B(n891), .A(n888), .S(n905), .Y(n895) );
  MUX2X1 U994 ( .B(n894), .A(n879), .S(n1001), .Y(n898) );
  MUX2X1 U995 ( .B(n897), .A(n834), .S(N24), .Y(n900) );
  INVX8 U996 ( .A(n908), .Y(n911) );
  INVX8 U997 ( .A(n908), .Y(n912) );
  INVX8 U998 ( .A(n908), .Y(n913) );
  INVX8 U999 ( .A(n916), .Y(n918) );
  INVX8 U1000 ( .A(n915), .Y(n919) );
  INVX8 U1001 ( .A(n915), .Y(n923) );
  INVX8 U1002 ( .A(n915), .Y(n924) );
  INVX8 U1003 ( .A(n915), .Y(n925) );
  INVX8 U1004 ( .A(n916), .Y(n926) );
  INVX8 U1005 ( .A(n915), .Y(n927) );
  INVX1 U1006 ( .A(N20), .Y(n1000) );
  INVX1 U1007 ( .A(N19), .Y(n999) );
  INVX1 U1008 ( .A(N18), .Y(n997) );
endmodule


module final_memory_3 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), err, .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<12> , \addr<11> , \addr<10> , \addr<9> , 
        \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , 
        \addr<2> , \addr<1> , \addr<0> }), wr, rd, enable, create_dump, 
    .bank_id({\bank_id<1> , \bank_id<0> }), clk, rst );
  input \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , \addr<12> , \addr<11> ,
         \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> , \addr<5> ,
         \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> , wr, rd, enable,
         create_dump, \bank_id<1> , \bank_id<0> , clk, rst;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , err;
  wire   n1046, rd0, wr0, rd1, wr1, \addr_1c<12> , \addr_1c<11> ,
         \addr_1c<10> , \addr_1c<9> , \addr_1c<8> , \addr_1c<7> , \addr_1c<6> ,
         \addr_1c<5> , \addr_1c<4> , \addr_1c<3> , \addr_1c<2> , \addr_1c<1> ,
         \addr_1c<0> , \data_in_1c<15> , \data_in_1c<14> , \data_in_1c<13> ,
         \data_in_1c<12> , \data_in_1c<11> , \data_in_1c<10> , \data_in_1c<9> ,
         \data_in_1c<8> , \data_in_1c<7> , \data_in_1c<6> , \data_in_1c<5> ,
         \data_in_1c<4> , \data_in_1c<3> , \data_in_1c<2> , \data_in_1c<1> ,
         \data_in_1c<0> , \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> ,
         \mem<0><3> , \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><7> ,
         \mem<1><6> , \mem<1><5> , \mem<1><4> , \mem<1><3> , \mem<1><2> ,
         \mem<1><1> , \mem<1><0> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><7> , \mem<3><6> , \mem<3><5> , \mem<3><4> , \mem<3><3> ,
         \mem<3><2> , \mem<3><1> , \mem<3><0> , \mem<4><7> , \mem<4><6> ,
         \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> , \mem<4><1> ,
         \mem<4><0> , \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> ,
         \mem<5><3> , \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><7> ,
         \mem<6><6> , \mem<6><5> , \mem<6><4> , \mem<6><3> , \mem<6><2> ,
         \mem<6><1> , \mem<6><0> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><7> , \mem<8><6> , \mem<8><5> , \mem<8><4> , \mem<8><3> ,
         \mem<8><2> , \mem<8><1> , \mem<8><0> , \mem<9><7> , \mem<9><6> ,
         \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> , \mem<9><1> ,
         \mem<9><0> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><7> ,
         \mem<11><6> , \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> ,
         \mem<11><1> , \mem<11><0> , \mem<12><7> , \mem<12><6> , \mem<12><5> ,
         \mem<12><4> , \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> ,
         \mem<13><7> , \mem<13><6> , \mem<13><5> , \mem<13><4> , \mem<13><3> ,
         \mem<13><2> , \mem<13><1> , \mem<13><0> , \mem<14><7> , \mem<14><6> ,
         \mem<14><5> , \mem<14><4> , \mem<14><3> , \mem<14><2> , \mem<14><1> ,
         \mem<14><0> , \mem<15><7> , \mem<15><6> , \mem<15><5> , \mem<15><4> ,
         \mem<15><3> , \mem<15><2> , \mem<15><1> , \mem<15><0> , \mem<16><7> ,
         \mem<16><6> , \mem<16><5> , \mem<16><4> , \mem<16><3> , \mem<16><2> ,
         \mem<16><1> , \mem<16><0> , \mem<17><7> , \mem<17><6> , \mem<17><5> ,
         \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> , \mem<17><0> ,
         \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> , \mem<18><3> ,
         \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><7> ,
         \mem<21><6> , \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> ,
         \mem<21><1> , \mem<21><0> , \mem<22><7> , \mem<22><6> , \mem<22><5> ,
         \mem<22><4> , \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> ,
         \mem<23><7> , \mem<23><6> , \mem<23><5> , \mem<23><4> , \mem<23><3> ,
         \mem<23><2> , \mem<23><1> , \mem<23><0> , \mem<24><7> , \mem<24><6> ,
         \mem<24><5> , \mem<24><4> , \mem<24><3> , \mem<24><2> , \mem<24><1> ,
         \mem<24><0> , \mem<25><7> , \mem<25><6> , \mem<25><5> , \mem<25><4> ,
         \mem<25><3> , \mem<25><2> , \mem<25><1> , \mem<25><0> , \mem<26><7> ,
         \mem<26><6> , \mem<26><5> , \mem<26><4> , \mem<26><3> , \mem<26><2> ,
         \mem<26><1> , \mem<26><0> , \mem<27><7> , \mem<27><6> , \mem<27><5> ,
         \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> , \mem<27><0> ,
         \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> , \mem<28><3> ,
         \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><7> ,
         \mem<31><6> , \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> ,
         \mem<31><1> , \mem<31><0> , \mem<32><7> , \mem<32><6> , \mem<32><5> ,
         \mem<32><4> , \mem<32><3> , \mem<32><2> , \mem<32><1> , \mem<32><0> ,
         \data_out_1c<15> , \data_out_1c<14> , \data_out_1c<13> ,
         \data_out_1c<12> , \data_out_1c<11> , \data_out_1c<10> ,
         \data_out_1c<9> , \data_out_1c<8> , rd2, wr2, rd3, wr3, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n373, n374, n375, n376, n377, n378, n380,
         n382, n383, n384, n385, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n403, n404, n405, n406, n407,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n584, n585, n586, n587,
         n588, n589, n590, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n50, n150, n189, n289, n348, n372, n379, n381, n386, n387,
         n401, n402, n409, n421, n422, n434, n435, n447, n448, n460, n461,
         n473, n474, n486, n487, n507, n508, n522, n523, n537, n538, n552,
         n553, n567, n568, n582, n583, n591, n592, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045;

  DFFPOSX1 \mem_reg<0><7>  ( .D(n870), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n869), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n868), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n867), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n866), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n865), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n864), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n863), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n862), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n861), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n860), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n859), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n858), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n857), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n856), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n855), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n854), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n853), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n852), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n851), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n850), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n849), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n848), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n847), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n846), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n845), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n844), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n843), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n842), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n841), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n840), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n839), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n838), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n837), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n836), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n835), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n834), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n833), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n832), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n831), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n830), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n829), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n828), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n827), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n826), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n825), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n824), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n823), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n822), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n821), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n820), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n819), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n818), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n817), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n816), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n815), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n814), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n813), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n812), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n811), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n810), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n809), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n808), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n807), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n806), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n805), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n804), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n803), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n802), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n801), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n800), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n799), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n798), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n797), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n796), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n795), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n794), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n793), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n792), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n791), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n790), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n789), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n788), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n787), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n786), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n785), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n784), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n783), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n782), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n781), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n780), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n779), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n778), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n777), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n776), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n775), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n774), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n773), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n772), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n771), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n770), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n769), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n768), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n767), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n766), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n765), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n764), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n763), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n762), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n761), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n760), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n759), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n758), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n757), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n756), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n755), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n754), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n753), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n752), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n751), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n750), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n749), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n748), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n747), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n746), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n745), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n744), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n743), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n742), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n741), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n740), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n739), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n738), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n737), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n736), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n735), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n734), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n733), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n732), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n731), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n730), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n729), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n728), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n727), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n726), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n725), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n724), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n723), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n722), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n721), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n720), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n719), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n718), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n717), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n716), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n715), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n714), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n713), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n712), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n711), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n710), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n709), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n708), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n707), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n706), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n705), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n704), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n703), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n702), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n701), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n700), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n699), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n698), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n697), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n696), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n695), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n694), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n693), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n692), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n691), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n690), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n689), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n688), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n687), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n686), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n685), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n684), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n683), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n682), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n681), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n680), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n679), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n678), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n677), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n676), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n675), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n674), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n673), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n672), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n671), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n670), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n669), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n668), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n667), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n666), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n665), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n664), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n663), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n662), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n661), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n660), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n659), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n658), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n657), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n656), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n655), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n654), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n653), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n652), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n651), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n650), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n649), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n648), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n647), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n646), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n645), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n644), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n643), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n642), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n641), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n640), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n639), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n638), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n637), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n636), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n635), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n634), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n633), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n632), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n631), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n630), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n629), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n628), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n627), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n626), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n625), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n624), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n623), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n622), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n621), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n620), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n619), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n618), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n617), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n616), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n615), .CLK(clk), .Q(\mem<31><0> ) );
  DFFPOSX1 \mem_reg<32><7>  ( .D(n614), .CLK(clk), .Q(\mem<32><7> ) );
  DFFPOSX1 \mem_reg<32><6>  ( .D(n613), .CLK(clk), .Q(\mem<32><6> ) );
  DFFPOSX1 \mem_reg<32><5>  ( .D(n612), .CLK(clk), .Q(\mem<32><5> ) );
  DFFPOSX1 \mem_reg<32><4>  ( .D(n611), .CLK(clk), .Q(\mem<32><4> ) );
  DFFPOSX1 \mem_reg<32><3>  ( .D(n610), .CLK(clk), .Q(\mem<32><3> ) );
  DFFPOSX1 \mem_reg<32><2>  ( .D(n609), .CLK(clk), .Q(\mem<32><2> ) );
  DFFPOSX1 \mem_reg<32><1>  ( .D(n608), .CLK(clk), .Q(\mem<32><1> ) );
  DFFPOSX1 \mem_reg<32><0>  ( .D(n607), .CLK(clk), .Q(\mem<32><0> ) );
  AND2X2 U9 ( .A(n413), .B(n414), .Y(n412) );
  AND2X2 U10 ( .A(n418), .B(n419), .Y(n417) );
  AND2X2 U11 ( .A(n426), .B(n427), .Y(n425) );
  AND2X2 U12 ( .A(n431), .B(n432), .Y(n430) );
  AND2X2 U13 ( .A(n439), .B(n440), .Y(n438) );
  AND2X2 U14 ( .A(n444), .B(n445), .Y(n443) );
  AND2X2 U15 ( .A(n452), .B(n453), .Y(n451) );
  AND2X2 U16 ( .A(n457), .B(n458), .Y(n456) );
  AND2X2 U17 ( .A(n465), .B(n466), .Y(n464) );
  AND2X2 U18 ( .A(n470), .B(n471), .Y(n469) );
  AND2X2 U19 ( .A(n478), .B(n479), .Y(n477) );
  AND2X2 U20 ( .A(n483), .B(n484), .Y(n482) );
  AND2X2 U21 ( .A(n491), .B(n492), .Y(n490) );
  AND2X2 U22 ( .A(n496), .B(n497), .Y(n495) );
  AND2X2 U30 ( .A(n588), .B(n1024), .Y(n248) );
  AND2X2 U31 ( .A(n589), .B(n1024), .Y(n91) );
  AND2X2 U32 ( .A(n588), .B(\addr_1c<0> ), .Y(n228) );
  AND2X2 U33 ( .A(n589), .B(\addr_1c<0> ), .Y(n71) );
  AND2X2 U34 ( .A(n596), .B(n597), .Y(n595) );
  AND2X2 U45 ( .A(n603), .B(n604), .Y(n602) );
  NOR3X1 U94 ( .A(n1044), .B(rd), .C(n963), .Y(wr0) );
  NOR3X1 U95 ( .A(n1045), .B(wr), .C(n963), .Y(rd0) );
  OAI21X1 U96 ( .A(n1011), .B(n1036), .C(n40), .Y(n607) );
  NAND2X1 U97 ( .A(\mem<32><0> ), .B(n1011), .Y(n40) );
  OAI21X1 U98 ( .A(n1011), .B(n1037), .C(n41), .Y(n608) );
  NAND2X1 U99 ( .A(\mem<32><1> ), .B(n1011), .Y(n41) );
  OAI21X1 U100 ( .A(n1011), .B(n1038), .C(n42), .Y(n609) );
  NAND2X1 U101 ( .A(\mem<32><2> ), .B(n1011), .Y(n42) );
  OAI21X1 U102 ( .A(n1011), .B(n1039), .C(n43), .Y(n610) );
  NAND2X1 U103 ( .A(\mem<32><3> ), .B(n1011), .Y(n43) );
  OAI21X1 U104 ( .A(n1011), .B(n1040), .C(n44), .Y(n611) );
  NAND2X1 U105 ( .A(\mem<32><4> ), .B(n1011), .Y(n44) );
  OAI21X1 U106 ( .A(n1011), .B(n1041), .C(n45), .Y(n612) );
  NAND2X1 U107 ( .A(\mem<32><5> ), .B(n1011), .Y(n45) );
  OAI21X1 U108 ( .A(n1011), .B(n1042), .C(n46), .Y(n613) );
  NAND2X1 U109 ( .A(\mem<32><6> ), .B(n1011), .Y(n46) );
  OAI21X1 U110 ( .A(n1011), .B(n1043), .C(n47), .Y(n614) );
  NAND2X1 U111 ( .A(\mem<32><7> ), .B(n1011), .Y(n47) );
  NAND3X1 U112 ( .A(n48), .B(n49), .C(n964), .Y(n39) );
  OAI21X1 U113 ( .A(n6), .B(n1028), .C(n51), .Y(n615) );
  NAND2X1 U114 ( .A(\mem<31><0> ), .B(n6), .Y(n51) );
  OAI21X1 U115 ( .A(n6), .B(n1029), .C(n52), .Y(n616) );
  NAND2X1 U116 ( .A(\mem<31><1> ), .B(n6), .Y(n52) );
  OAI21X1 U117 ( .A(n6), .B(n1030), .C(n53), .Y(n617) );
  NAND2X1 U118 ( .A(\mem<31><2> ), .B(n6), .Y(n53) );
  OAI21X1 U119 ( .A(n6), .B(n1031), .C(n54), .Y(n618) );
  NAND2X1 U120 ( .A(\mem<31><3> ), .B(n6), .Y(n54) );
  OAI21X1 U121 ( .A(n6), .B(n1032), .C(n55), .Y(n619) );
  NAND2X1 U122 ( .A(\mem<31><4> ), .B(n6), .Y(n55) );
  OAI21X1 U123 ( .A(n6), .B(n1033), .C(n56), .Y(n620) );
  NAND2X1 U124 ( .A(\mem<31><5> ), .B(n6), .Y(n56) );
  OAI21X1 U125 ( .A(n6), .B(n1034), .C(n57), .Y(n621) );
  NAND2X1 U126 ( .A(\mem<31><6> ), .B(n6), .Y(n57) );
  OAI21X1 U127 ( .A(n6), .B(n1035), .C(n58), .Y(n622) );
  NAND2X1 U128 ( .A(\mem<31><7> ), .B(n6), .Y(n58) );
  OAI21X1 U130 ( .A(n1036), .B(n1010), .C(n62), .Y(n623) );
  NAND2X1 U131 ( .A(\mem<30><0> ), .B(n1010), .Y(n62) );
  OAI21X1 U132 ( .A(n1037), .B(n1009), .C(n63), .Y(n624) );
  NAND2X1 U133 ( .A(\mem<30><1> ), .B(n1010), .Y(n63) );
  OAI21X1 U134 ( .A(n1038), .B(n1009), .C(n64), .Y(n625) );
  NAND2X1 U135 ( .A(\mem<30><2> ), .B(n1010), .Y(n64) );
  OAI21X1 U136 ( .A(n1039), .B(n1009), .C(n65), .Y(n626) );
  NAND2X1 U137 ( .A(\mem<30><3> ), .B(n1010), .Y(n65) );
  OAI21X1 U138 ( .A(n1040), .B(n1009), .C(n66), .Y(n627) );
  NAND2X1 U139 ( .A(\mem<30><4> ), .B(n1010), .Y(n66) );
  OAI21X1 U140 ( .A(n1041), .B(n1009), .C(n67), .Y(n628) );
  NAND2X1 U141 ( .A(\mem<30><5> ), .B(n1010), .Y(n67) );
  OAI21X1 U142 ( .A(n1042), .B(n1009), .C(n68), .Y(n629) );
  NAND2X1 U143 ( .A(\mem<30><6> ), .B(n1010), .Y(n68) );
  OAI21X1 U144 ( .A(n1043), .B(n1009), .C(n69), .Y(n630) );
  NAND2X1 U145 ( .A(\mem<30><7> ), .B(n1010), .Y(n69) );
  NAND3X1 U146 ( .A(n70), .B(n48), .C(n71), .Y(n61) );
  OAI21X1 U147 ( .A(n1028), .B(n1008), .C(n73), .Y(n631) );
  NAND2X1 U148 ( .A(\mem<29><0> ), .B(n1008), .Y(n73) );
  OAI21X1 U149 ( .A(n1029), .B(n1008), .C(n74), .Y(n632) );
  NAND2X1 U150 ( .A(\mem<29><1> ), .B(n1008), .Y(n74) );
  OAI21X1 U151 ( .A(n1030), .B(n1008), .C(n75), .Y(n633) );
  NAND2X1 U152 ( .A(\mem<29><2> ), .B(n1008), .Y(n75) );
  OAI21X1 U153 ( .A(n1031), .B(n1008), .C(n76), .Y(n634) );
  NAND2X1 U154 ( .A(\mem<29><3> ), .B(n1008), .Y(n76) );
  OAI21X1 U155 ( .A(n1032), .B(n1008), .C(n77), .Y(n635) );
  NAND2X1 U156 ( .A(\mem<29><4> ), .B(n1008), .Y(n77) );
  OAI21X1 U157 ( .A(n1033), .B(n1008), .C(n78), .Y(n636) );
  NAND2X1 U158 ( .A(\mem<29><5> ), .B(n1008), .Y(n78) );
  OAI21X1 U159 ( .A(n1034), .B(n1008), .C(n79), .Y(n637) );
  NAND2X1 U160 ( .A(\mem<29><6> ), .B(n1008), .Y(n79) );
  OAI21X1 U161 ( .A(n1035), .B(n1008), .C(n80), .Y(n638) );
  NAND2X1 U162 ( .A(\mem<29><7> ), .B(n1008), .Y(n80) );
  NAND3X1 U163 ( .A(n973), .B(n48), .C(n81), .Y(n72) );
  OAI21X1 U164 ( .A(n1036), .B(n1007), .C(n83), .Y(n639) );
  NAND2X1 U165 ( .A(\mem<28><0> ), .B(n1007), .Y(n83) );
  OAI21X1 U166 ( .A(n1037), .B(n1006), .C(n84), .Y(n640) );
  NAND2X1 U167 ( .A(\mem<28><1> ), .B(n1007), .Y(n84) );
  OAI21X1 U168 ( .A(n1038), .B(n1006), .C(n85), .Y(n641) );
  NAND2X1 U169 ( .A(\mem<28><2> ), .B(n1007), .Y(n85) );
  OAI21X1 U170 ( .A(n1039), .B(n1006), .C(n86), .Y(n642) );
  NAND2X1 U171 ( .A(\mem<28><3> ), .B(n1007), .Y(n86) );
  OAI21X1 U172 ( .A(n1040), .B(n1006), .C(n87), .Y(n643) );
  NAND2X1 U173 ( .A(\mem<28><4> ), .B(n1007), .Y(n87) );
  OAI21X1 U174 ( .A(n1041), .B(n1006), .C(n88), .Y(n644) );
  NAND2X1 U175 ( .A(\mem<28><5> ), .B(n1007), .Y(n88) );
  OAI21X1 U176 ( .A(n1042), .B(n1006), .C(n89), .Y(n645) );
  NAND2X1 U177 ( .A(\mem<28><6> ), .B(n1007), .Y(n89) );
  OAI21X1 U178 ( .A(n1043), .B(n1006), .C(n90), .Y(n646) );
  NAND2X1 U179 ( .A(\mem<28><7> ), .B(n1007), .Y(n90) );
  NAND3X1 U180 ( .A(n70), .B(n48), .C(n91), .Y(n82) );
  OAI21X1 U181 ( .A(n1028), .B(n1005), .C(n93), .Y(n647) );
  NAND2X1 U182 ( .A(\mem<27><0> ), .B(n1005), .Y(n93) );
  OAI21X1 U183 ( .A(n1029), .B(n1005), .C(n94), .Y(n648) );
  NAND2X1 U184 ( .A(\mem<27><1> ), .B(n1005), .Y(n94) );
  OAI21X1 U185 ( .A(n1030), .B(n1005), .C(n95), .Y(n649) );
  NAND2X1 U186 ( .A(\mem<27><2> ), .B(n1005), .Y(n95) );
  OAI21X1 U187 ( .A(n1031), .B(n1005), .C(n96), .Y(n650) );
  NAND2X1 U188 ( .A(\mem<27><3> ), .B(n1005), .Y(n96) );
  OAI21X1 U189 ( .A(n1032), .B(n1005), .C(n97), .Y(n651) );
  NAND2X1 U190 ( .A(\mem<27><4> ), .B(n1005), .Y(n97) );
  OAI21X1 U191 ( .A(n1033), .B(n1005), .C(n98), .Y(n652) );
  NAND2X1 U192 ( .A(\mem<27><5> ), .B(n1005), .Y(n98) );
  OAI21X1 U193 ( .A(n1034), .B(n1005), .C(n99), .Y(n653) );
  NAND2X1 U194 ( .A(\mem<27><6> ), .B(n1005), .Y(n99) );
  OAI21X1 U195 ( .A(n1035), .B(n1005), .C(n100), .Y(n654) );
  NAND2X1 U196 ( .A(\mem<27><7> ), .B(n1005), .Y(n100) );
  NAND3X1 U197 ( .A(n973), .B(n48), .C(n101), .Y(n92) );
  OAI21X1 U198 ( .A(n1036), .B(n1004), .C(n103), .Y(n655) );
  NAND2X1 U199 ( .A(\mem<26><0> ), .B(n1004), .Y(n103) );
  OAI21X1 U200 ( .A(n1037), .B(n1003), .C(n104), .Y(n656) );
  NAND2X1 U201 ( .A(\mem<26><1> ), .B(n1004), .Y(n104) );
  OAI21X1 U202 ( .A(n1038), .B(n1003), .C(n105), .Y(n657) );
  NAND2X1 U203 ( .A(\mem<26><2> ), .B(n1004), .Y(n105) );
  OAI21X1 U204 ( .A(n1039), .B(n1003), .C(n106), .Y(n658) );
  NAND2X1 U205 ( .A(\mem<26><3> ), .B(n1004), .Y(n106) );
  OAI21X1 U206 ( .A(n1040), .B(n1003), .C(n107), .Y(n659) );
  NAND2X1 U207 ( .A(\mem<26><4> ), .B(n1004), .Y(n107) );
  OAI21X1 U208 ( .A(n1041), .B(n1003), .C(n108), .Y(n660) );
  NAND2X1 U209 ( .A(\mem<26><5> ), .B(n1004), .Y(n108) );
  OAI21X1 U210 ( .A(n1042), .B(n1003), .C(n109), .Y(n661) );
  NAND2X1 U211 ( .A(\mem<26><6> ), .B(n1004), .Y(n109) );
  OAI21X1 U212 ( .A(n1043), .B(n1003), .C(n110), .Y(n662) );
  NAND2X1 U213 ( .A(\mem<26><7> ), .B(n1004), .Y(n110) );
  NAND3X1 U214 ( .A(n71), .B(n48), .C(n111), .Y(n102) );
  OAI21X1 U215 ( .A(n1028), .B(n1002), .C(n113), .Y(n663) );
  NAND2X1 U216 ( .A(\mem<25><0> ), .B(n1002), .Y(n113) );
  OAI21X1 U217 ( .A(n1029), .B(n1002), .C(n114), .Y(n664) );
  NAND2X1 U218 ( .A(\mem<25><1> ), .B(n1002), .Y(n114) );
  OAI21X1 U219 ( .A(n1030), .B(n1002), .C(n115), .Y(n665) );
  NAND2X1 U220 ( .A(\mem<25><2> ), .B(n1002), .Y(n115) );
  OAI21X1 U221 ( .A(n1031), .B(n1002), .C(n116), .Y(n666) );
  NAND2X1 U222 ( .A(\mem<25><3> ), .B(n1002), .Y(n116) );
  OAI21X1 U223 ( .A(n1032), .B(n1002), .C(n117), .Y(n667) );
  NAND2X1 U224 ( .A(\mem<25><4> ), .B(n1002), .Y(n117) );
  OAI21X1 U225 ( .A(n1033), .B(n1002), .C(n118), .Y(n668) );
  NAND2X1 U226 ( .A(\mem<25><5> ), .B(n1002), .Y(n118) );
  OAI21X1 U227 ( .A(n1034), .B(n1002), .C(n119), .Y(n669) );
  NAND2X1 U228 ( .A(\mem<25><6> ), .B(n1002), .Y(n119) );
  OAI21X1 U229 ( .A(n1035), .B(n1002), .C(n120), .Y(n670) );
  NAND2X1 U230 ( .A(\mem<25><7> ), .B(n1002), .Y(n120) );
  NAND3X1 U231 ( .A(n973), .B(n48), .C(n121), .Y(n112) );
  OAI21X1 U232 ( .A(n1036), .B(n1001), .C(n123), .Y(n671) );
  NAND2X1 U233 ( .A(\mem<24><0> ), .B(n1001), .Y(n123) );
  OAI21X1 U234 ( .A(n1037), .B(n1000), .C(n124), .Y(n672) );
  NAND2X1 U235 ( .A(\mem<24><1> ), .B(n1001), .Y(n124) );
  OAI21X1 U236 ( .A(n1038), .B(n1000), .C(n125), .Y(n673) );
  NAND2X1 U237 ( .A(\mem<24><2> ), .B(n1001), .Y(n125) );
  OAI21X1 U238 ( .A(n1039), .B(n1000), .C(n126), .Y(n674) );
  NAND2X1 U239 ( .A(\mem<24><3> ), .B(n1001), .Y(n126) );
  OAI21X1 U240 ( .A(n1040), .B(n1000), .C(n127), .Y(n675) );
  NAND2X1 U241 ( .A(\mem<24><4> ), .B(n1001), .Y(n127) );
  OAI21X1 U242 ( .A(n1041), .B(n1000), .C(n128), .Y(n676) );
  NAND2X1 U243 ( .A(\mem<24><5> ), .B(n1001), .Y(n128) );
  OAI21X1 U244 ( .A(n1042), .B(n1000), .C(n129), .Y(n677) );
  NAND2X1 U245 ( .A(\mem<24><6> ), .B(n1001), .Y(n129) );
  OAI21X1 U246 ( .A(n1043), .B(n1000), .C(n130), .Y(n678) );
  NAND2X1 U247 ( .A(\mem<24><7> ), .B(n1001), .Y(n130) );
  NAND3X1 U248 ( .A(n91), .B(n48), .C(n111), .Y(n122) );
  OAI21X1 U249 ( .A(n1028), .B(n999), .C(n132), .Y(n679) );
  NAND2X1 U250 ( .A(\mem<23><0> ), .B(n999), .Y(n132) );
  OAI21X1 U251 ( .A(n1029), .B(n999), .C(n133), .Y(n680) );
  NAND2X1 U252 ( .A(\mem<23><1> ), .B(n999), .Y(n133) );
  OAI21X1 U253 ( .A(n1030), .B(n999), .C(n134), .Y(n681) );
  NAND2X1 U254 ( .A(\mem<23><2> ), .B(n999), .Y(n134) );
  OAI21X1 U255 ( .A(n1031), .B(n999), .C(n135), .Y(n682) );
  NAND2X1 U256 ( .A(\mem<23><3> ), .B(n999), .Y(n135) );
  OAI21X1 U257 ( .A(n1032), .B(n999), .C(n136), .Y(n683) );
  NAND2X1 U258 ( .A(\mem<23><4> ), .B(n999), .Y(n136) );
  OAI21X1 U259 ( .A(n1033), .B(n999), .C(n137), .Y(n684) );
  NAND2X1 U260 ( .A(\mem<23><5> ), .B(n999), .Y(n137) );
  OAI21X1 U261 ( .A(n1034), .B(n999), .C(n138), .Y(n685) );
  NAND2X1 U262 ( .A(\mem<23><6> ), .B(n999), .Y(n138) );
  OAI21X1 U263 ( .A(n1035), .B(n999), .C(n139), .Y(n686) );
  NAND2X1 U264 ( .A(\mem<23><7> ), .B(n999), .Y(n139) );
  NAND3X1 U265 ( .A(n973), .B(n48), .C(n140), .Y(n131) );
  OAI21X1 U266 ( .A(n1036), .B(n998), .C(n142), .Y(n687) );
  NAND2X1 U267 ( .A(\mem<22><0> ), .B(n998), .Y(n142) );
  OAI21X1 U268 ( .A(n1037), .B(n998), .C(n143), .Y(n688) );
  NAND2X1 U269 ( .A(\mem<22><1> ), .B(n998), .Y(n143) );
  OAI21X1 U270 ( .A(n1038), .B(n998), .C(n144), .Y(n689) );
  NAND2X1 U271 ( .A(\mem<22><2> ), .B(n998), .Y(n144) );
  OAI21X1 U272 ( .A(n1039), .B(n998), .C(n145), .Y(n690) );
  NAND2X1 U273 ( .A(\mem<22><3> ), .B(n998), .Y(n145) );
  OAI21X1 U274 ( .A(n1040), .B(n998), .C(n146), .Y(n691) );
  NAND2X1 U275 ( .A(\mem<22><4> ), .B(n998), .Y(n146) );
  OAI21X1 U276 ( .A(n1041), .B(n998), .C(n147), .Y(n692) );
  NAND2X1 U277 ( .A(\mem<22><5> ), .B(n998), .Y(n147) );
  OAI21X1 U278 ( .A(n1042), .B(n998), .C(n148), .Y(n693) );
  NAND2X1 U279 ( .A(\mem<22><6> ), .B(n998), .Y(n148) );
  OAI21X1 U280 ( .A(n1043), .B(n998), .C(n149), .Y(n694) );
  NAND2X1 U281 ( .A(\mem<22><7> ), .B(n998), .Y(n149) );
  NAND3X1 U282 ( .A(n71), .B(n48), .C(n969), .Y(n141) );
  OAI21X1 U283 ( .A(n1028), .B(n997), .C(n152), .Y(n695) );
  NAND2X1 U284 ( .A(\mem<21><0> ), .B(n997), .Y(n152) );
  OAI21X1 U285 ( .A(n1029), .B(n997), .C(n153), .Y(n696) );
  NAND2X1 U286 ( .A(\mem<21><1> ), .B(n997), .Y(n153) );
  OAI21X1 U287 ( .A(n1030), .B(n997), .C(n154), .Y(n697) );
  NAND2X1 U288 ( .A(\mem<21><2> ), .B(n997), .Y(n154) );
  OAI21X1 U289 ( .A(n1031), .B(n997), .C(n155), .Y(n698) );
  NAND2X1 U290 ( .A(\mem<21><3> ), .B(n997), .Y(n155) );
  OAI21X1 U291 ( .A(n1032), .B(n997), .C(n156), .Y(n699) );
  NAND2X1 U292 ( .A(\mem<21><4> ), .B(n997), .Y(n156) );
  OAI21X1 U293 ( .A(n1033), .B(n997), .C(n157), .Y(n700) );
  NAND2X1 U294 ( .A(\mem<21><5> ), .B(n997), .Y(n157) );
  OAI21X1 U295 ( .A(n1034), .B(n997), .C(n158), .Y(n701) );
  NAND2X1 U296 ( .A(\mem<21><6> ), .B(n997), .Y(n158) );
  OAI21X1 U297 ( .A(n1035), .B(n997), .C(n159), .Y(n702) );
  NAND2X1 U298 ( .A(\mem<21><7> ), .B(n997), .Y(n159) );
  NAND3X1 U299 ( .A(n973), .B(n48), .C(n160), .Y(n151) );
  OAI21X1 U300 ( .A(n1036), .B(n996), .C(n162), .Y(n703) );
  NAND2X1 U301 ( .A(\mem<20><0> ), .B(n996), .Y(n162) );
  OAI21X1 U302 ( .A(n1037), .B(n996), .C(n163), .Y(n704) );
  NAND2X1 U303 ( .A(\mem<20><1> ), .B(n996), .Y(n163) );
  OAI21X1 U304 ( .A(n1038), .B(n996), .C(n164), .Y(n705) );
  NAND2X1 U305 ( .A(\mem<20><2> ), .B(n996), .Y(n164) );
  OAI21X1 U306 ( .A(n1039), .B(n996), .C(n165), .Y(n706) );
  NAND2X1 U307 ( .A(\mem<20><3> ), .B(n996), .Y(n165) );
  OAI21X1 U308 ( .A(n1040), .B(n996), .C(n166), .Y(n707) );
  NAND2X1 U309 ( .A(\mem<20><4> ), .B(n996), .Y(n166) );
  OAI21X1 U310 ( .A(n1041), .B(n996), .C(n167), .Y(n708) );
  NAND2X1 U311 ( .A(\mem<20><5> ), .B(n996), .Y(n167) );
  OAI21X1 U312 ( .A(n1042), .B(n996), .C(n168), .Y(n709) );
  NAND2X1 U313 ( .A(\mem<20><6> ), .B(n996), .Y(n168) );
  OAI21X1 U314 ( .A(n1043), .B(n996), .C(n169), .Y(n710) );
  NAND2X1 U315 ( .A(\mem<20><7> ), .B(n996), .Y(n169) );
  NAND3X1 U316 ( .A(n91), .B(n48), .C(n969), .Y(n161) );
  OAI21X1 U317 ( .A(n1028), .B(n995), .C(n171), .Y(n711) );
  NAND2X1 U318 ( .A(\mem<19><0> ), .B(n995), .Y(n171) );
  OAI21X1 U319 ( .A(n1029), .B(n995), .C(n172), .Y(n712) );
  NAND2X1 U320 ( .A(\mem<19><1> ), .B(n995), .Y(n172) );
  OAI21X1 U321 ( .A(n1030), .B(n995), .C(n173), .Y(n713) );
  NAND2X1 U322 ( .A(\mem<19><2> ), .B(n995), .Y(n173) );
  OAI21X1 U323 ( .A(n1031), .B(n995), .C(n174), .Y(n714) );
  NAND2X1 U324 ( .A(\mem<19><3> ), .B(n995), .Y(n174) );
  OAI21X1 U325 ( .A(n1032), .B(n995), .C(n175), .Y(n715) );
  NAND2X1 U326 ( .A(\mem<19><4> ), .B(n995), .Y(n175) );
  OAI21X1 U327 ( .A(n1033), .B(n995), .C(n176), .Y(n716) );
  NAND2X1 U328 ( .A(\mem<19><5> ), .B(n995), .Y(n176) );
  OAI21X1 U329 ( .A(n1034), .B(n995), .C(n177), .Y(n717) );
  NAND2X1 U330 ( .A(\mem<19><6> ), .B(n995), .Y(n177) );
  OAI21X1 U331 ( .A(n1035), .B(n995), .C(n178), .Y(n718) );
  NAND2X1 U332 ( .A(\mem<19><7> ), .B(n995), .Y(n178) );
  NAND3X1 U333 ( .A(n973), .B(n48), .C(n179), .Y(n170) );
  OAI21X1 U334 ( .A(n1036), .B(n994), .C(n181), .Y(n719) );
  NAND2X1 U335 ( .A(\mem<18><0> ), .B(n994), .Y(n181) );
  OAI21X1 U336 ( .A(n1037), .B(n994), .C(n182), .Y(n720) );
  NAND2X1 U337 ( .A(\mem<18><1> ), .B(n994), .Y(n182) );
  OAI21X1 U338 ( .A(n1038), .B(n994), .C(n183), .Y(n721) );
  NAND2X1 U339 ( .A(\mem<18><2> ), .B(n994), .Y(n183) );
  OAI21X1 U340 ( .A(n1039), .B(n994), .C(n184), .Y(n722) );
  NAND2X1 U341 ( .A(\mem<18><3> ), .B(n994), .Y(n184) );
  OAI21X1 U342 ( .A(n1040), .B(n994), .C(n185), .Y(n723) );
  NAND2X1 U343 ( .A(\mem<18><4> ), .B(n994), .Y(n185) );
  OAI21X1 U344 ( .A(n1041), .B(n994), .C(n186), .Y(n724) );
  NAND2X1 U345 ( .A(\mem<18><5> ), .B(n994), .Y(n186) );
  OAI21X1 U346 ( .A(n1042), .B(n994), .C(n187), .Y(n725) );
  NAND2X1 U347 ( .A(\mem<18><6> ), .B(n994), .Y(n187) );
  OAI21X1 U348 ( .A(n1043), .B(n994), .C(n188), .Y(n726) );
  NAND2X1 U349 ( .A(\mem<18><7> ), .B(n994), .Y(n188) );
  NAND3X1 U350 ( .A(n71), .B(n48), .C(n967), .Y(n180) );
  OAI21X1 U351 ( .A(n1028), .B(n993), .C(n191), .Y(n727) );
  NAND2X1 U352 ( .A(\mem<17><0> ), .B(n993), .Y(n191) );
  OAI21X1 U353 ( .A(n1029), .B(n993), .C(n192), .Y(n728) );
  NAND2X1 U354 ( .A(\mem<17><1> ), .B(n993), .Y(n192) );
  OAI21X1 U355 ( .A(n1030), .B(n993), .C(n193), .Y(n729) );
  NAND2X1 U356 ( .A(\mem<17><2> ), .B(n993), .Y(n193) );
  OAI21X1 U357 ( .A(n1031), .B(n993), .C(n194), .Y(n730) );
  NAND2X1 U358 ( .A(\mem<17><3> ), .B(n993), .Y(n194) );
  OAI21X1 U359 ( .A(n1032), .B(n993), .C(n195), .Y(n731) );
  NAND2X1 U360 ( .A(\mem<17><4> ), .B(n993), .Y(n195) );
  OAI21X1 U361 ( .A(n1033), .B(n993), .C(n196), .Y(n732) );
  NAND2X1 U362 ( .A(\mem<17><5> ), .B(n993), .Y(n196) );
  OAI21X1 U363 ( .A(n1034), .B(n993), .C(n197), .Y(n733) );
  NAND2X1 U364 ( .A(\mem<17><6> ), .B(n993), .Y(n197) );
  OAI21X1 U365 ( .A(n1035), .B(n993), .C(n198), .Y(n734) );
  NAND2X1 U366 ( .A(\mem<17><7> ), .B(n993), .Y(n198) );
  NAND3X1 U367 ( .A(n973), .B(n48), .C(n199), .Y(n190) );
  OAI21X1 U368 ( .A(n1036), .B(n992), .C(n201), .Y(n735) );
  NAND2X1 U369 ( .A(\mem<16><0> ), .B(n992), .Y(n201) );
  OAI21X1 U370 ( .A(n1037), .B(n992), .C(n202), .Y(n736) );
  NAND2X1 U371 ( .A(\mem<16><1> ), .B(n992), .Y(n202) );
  OAI21X1 U372 ( .A(n1038), .B(n992), .C(n203), .Y(n737) );
  NAND2X1 U373 ( .A(\mem<16><2> ), .B(n992), .Y(n203) );
  OAI21X1 U374 ( .A(n1039), .B(n992), .C(n204), .Y(n738) );
  NAND2X1 U375 ( .A(\mem<16><3> ), .B(n992), .Y(n204) );
  OAI21X1 U376 ( .A(n1040), .B(n992), .C(n205), .Y(n739) );
  NAND2X1 U377 ( .A(\mem<16><4> ), .B(n992), .Y(n205) );
  OAI21X1 U378 ( .A(n1041), .B(n992), .C(n206), .Y(n740) );
  NAND2X1 U379 ( .A(\mem<16><5> ), .B(n992), .Y(n206) );
  OAI21X1 U380 ( .A(n1042), .B(n992), .C(n207), .Y(n741) );
  NAND2X1 U381 ( .A(\mem<16><6> ), .B(n992), .Y(n207) );
  OAI21X1 U382 ( .A(n1043), .B(n992), .C(n208), .Y(n742) );
  NAND2X1 U383 ( .A(\mem<16><7> ), .B(n992), .Y(n208) );
  NAND3X1 U384 ( .A(n91), .B(n48), .C(n967), .Y(n200) );
  OAI21X1 U385 ( .A(n1028), .B(n991), .C(n210), .Y(n743) );
  NAND2X1 U386 ( .A(\mem<15><0> ), .B(n991), .Y(n210) );
  OAI21X1 U387 ( .A(n1029), .B(n991), .C(n211), .Y(n744) );
  NAND2X1 U388 ( .A(\mem<15><1> ), .B(n991), .Y(n211) );
  OAI21X1 U389 ( .A(n1030), .B(n991), .C(n212), .Y(n745) );
  NAND2X1 U390 ( .A(\mem<15><2> ), .B(n991), .Y(n212) );
  OAI21X1 U391 ( .A(n1031), .B(n991), .C(n213), .Y(n746) );
  NAND2X1 U392 ( .A(\mem<15><3> ), .B(n991), .Y(n213) );
  OAI21X1 U393 ( .A(n1032), .B(n991), .C(n214), .Y(n747) );
  NAND2X1 U394 ( .A(\mem<15><4> ), .B(n991), .Y(n214) );
  OAI21X1 U395 ( .A(n1033), .B(n991), .C(n215), .Y(n748) );
  NAND2X1 U396 ( .A(\mem<15><5> ), .B(n991), .Y(n215) );
  OAI21X1 U397 ( .A(n1034), .B(n991), .C(n216), .Y(n749) );
  NAND2X1 U398 ( .A(\mem<15><6> ), .B(n991), .Y(n216) );
  OAI21X1 U399 ( .A(n1035), .B(n991), .C(n217), .Y(n750) );
  NAND2X1 U400 ( .A(\mem<15><7> ), .B(n991), .Y(n217) );
  NAND3X1 U401 ( .A(n973), .B(n48), .C(n218), .Y(n209) );
  OAI21X1 U402 ( .A(n1036), .B(n990), .C(n220), .Y(n751) );
  NAND2X1 U403 ( .A(\mem<14><0> ), .B(n990), .Y(n220) );
  OAI21X1 U404 ( .A(n1037), .B(n989), .C(n221), .Y(n752) );
  NAND2X1 U405 ( .A(\mem<14><1> ), .B(n990), .Y(n221) );
  OAI21X1 U406 ( .A(n1038), .B(n989), .C(n222), .Y(n753) );
  NAND2X1 U407 ( .A(\mem<14><2> ), .B(n990), .Y(n222) );
  OAI21X1 U408 ( .A(n1039), .B(n989), .C(n223), .Y(n754) );
  NAND2X1 U409 ( .A(\mem<14><3> ), .B(n990), .Y(n223) );
  OAI21X1 U410 ( .A(n1040), .B(n989), .C(n224), .Y(n755) );
  NAND2X1 U411 ( .A(\mem<14><4> ), .B(n990), .Y(n224) );
  OAI21X1 U412 ( .A(n1041), .B(n989), .C(n225), .Y(n756) );
  NAND2X1 U413 ( .A(\mem<14><5> ), .B(n990), .Y(n225) );
  OAI21X1 U414 ( .A(n1042), .B(n989), .C(n226), .Y(n757) );
  NAND2X1 U415 ( .A(\mem<14><6> ), .B(n990), .Y(n226) );
  OAI21X1 U416 ( .A(n1043), .B(n989), .C(n227), .Y(n758) );
  NAND2X1 U417 ( .A(\mem<14><7> ), .B(n990), .Y(n227) );
  NAND3X1 U418 ( .A(n70), .B(n48), .C(n228), .Y(n219) );
  OAI21X1 U419 ( .A(n1028), .B(n988), .C(n230), .Y(n759) );
  NAND2X1 U420 ( .A(\mem<13><0> ), .B(n988), .Y(n230) );
  OAI21X1 U421 ( .A(n1029), .B(n988), .C(n231), .Y(n760) );
  NAND2X1 U422 ( .A(\mem<13><1> ), .B(n988), .Y(n231) );
  OAI21X1 U423 ( .A(n1030), .B(n988), .C(n232), .Y(n761) );
  NAND2X1 U424 ( .A(\mem<13><2> ), .B(n988), .Y(n232) );
  OAI21X1 U425 ( .A(n1031), .B(n988), .C(n233), .Y(n762) );
  NAND2X1 U426 ( .A(\mem<13><3> ), .B(n988), .Y(n233) );
  OAI21X1 U427 ( .A(n1032), .B(n988), .C(n234), .Y(n763) );
  NAND2X1 U428 ( .A(\mem<13><4> ), .B(n988), .Y(n234) );
  OAI21X1 U429 ( .A(n1033), .B(n988), .C(n235), .Y(n764) );
  NAND2X1 U430 ( .A(\mem<13><5> ), .B(n988), .Y(n235) );
  OAI21X1 U431 ( .A(n1034), .B(n988), .C(n236), .Y(n765) );
  NAND2X1 U432 ( .A(\mem<13><6> ), .B(n988), .Y(n236) );
  OAI21X1 U433 ( .A(n1035), .B(n988), .C(n237), .Y(n766) );
  NAND2X1 U434 ( .A(\mem<13><7> ), .B(n988), .Y(n237) );
  NAND3X1 U435 ( .A(n973), .B(n48), .C(n238), .Y(n229) );
  OAI21X1 U436 ( .A(n1036), .B(n987), .C(n240), .Y(n767) );
  NAND2X1 U437 ( .A(\mem<12><0> ), .B(n987), .Y(n240) );
  OAI21X1 U438 ( .A(n1037), .B(n986), .C(n241), .Y(n768) );
  NAND2X1 U439 ( .A(\mem<12><1> ), .B(n987), .Y(n241) );
  OAI21X1 U440 ( .A(n1038), .B(n986), .C(n242), .Y(n769) );
  NAND2X1 U441 ( .A(\mem<12><2> ), .B(n987), .Y(n242) );
  OAI21X1 U442 ( .A(n1039), .B(n986), .C(n243), .Y(n770) );
  NAND2X1 U443 ( .A(\mem<12><3> ), .B(n987), .Y(n243) );
  OAI21X1 U444 ( .A(n1040), .B(n986), .C(n244), .Y(n771) );
  NAND2X1 U445 ( .A(\mem<12><4> ), .B(n987), .Y(n244) );
  OAI21X1 U446 ( .A(n1041), .B(n986), .C(n245), .Y(n772) );
  NAND2X1 U447 ( .A(\mem<12><5> ), .B(n987), .Y(n245) );
  OAI21X1 U448 ( .A(n1042), .B(n986), .C(n246), .Y(n773) );
  NAND2X1 U449 ( .A(\mem<12><6> ), .B(n987), .Y(n246) );
  OAI21X1 U450 ( .A(n1043), .B(n986), .C(n247), .Y(n774) );
  NAND2X1 U451 ( .A(\mem<12><7> ), .B(n987), .Y(n247) );
  NAND3X1 U452 ( .A(n70), .B(n48), .C(n248), .Y(n239) );
  OAI21X1 U453 ( .A(n1028), .B(n985), .C(n251), .Y(n775) );
  NAND2X1 U454 ( .A(\mem<11><0> ), .B(n985), .Y(n251) );
  OAI21X1 U455 ( .A(n1029), .B(n985), .C(n252), .Y(n776) );
  NAND2X1 U456 ( .A(\mem<11><1> ), .B(n985), .Y(n252) );
  OAI21X1 U457 ( .A(n1030), .B(n985), .C(n253), .Y(n777) );
  NAND2X1 U458 ( .A(\mem<11><2> ), .B(n985), .Y(n253) );
  OAI21X1 U459 ( .A(n1031), .B(n985), .C(n254), .Y(n778) );
  NAND2X1 U460 ( .A(\mem<11><3> ), .B(n985), .Y(n254) );
  OAI21X1 U461 ( .A(n1032), .B(n985), .C(n255), .Y(n779) );
  NAND2X1 U462 ( .A(\mem<11><4> ), .B(n985), .Y(n255) );
  OAI21X1 U463 ( .A(n1033), .B(n985), .C(n256), .Y(n780) );
  NAND2X1 U464 ( .A(\mem<11><5> ), .B(n985), .Y(n256) );
  OAI21X1 U465 ( .A(n1034), .B(n985), .C(n257), .Y(n781) );
  NAND2X1 U466 ( .A(\mem<11><6> ), .B(n985), .Y(n257) );
  OAI21X1 U467 ( .A(n1035), .B(n985), .C(n258), .Y(n782) );
  NAND2X1 U468 ( .A(\mem<11><7> ), .B(n985), .Y(n258) );
  NAND3X1 U469 ( .A(n973), .B(n48), .C(n259), .Y(n250) );
  OAI21X1 U470 ( .A(n1036), .B(n984), .C(n261), .Y(n783) );
  NAND2X1 U471 ( .A(\mem<10><0> ), .B(n984), .Y(n261) );
  OAI21X1 U472 ( .A(n1037), .B(n983), .C(n262), .Y(n784) );
  NAND2X1 U473 ( .A(\mem<10><1> ), .B(n984), .Y(n262) );
  OAI21X1 U474 ( .A(n1038), .B(n983), .C(n263), .Y(n785) );
  NAND2X1 U475 ( .A(\mem<10><2> ), .B(n984), .Y(n263) );
  OAI21X1 U476 ( .A(n1039), .B(n983), .C(n264), .Y(n786) );
  NAND2X1 U477 ( .A(\mem<10><3> ), .B(n984), .Y(n264) );
  OAI21X1 U478 ( .A(n1040), .B(n983), .C(n265), .Y(n787) );
  NAND2X1 U479 ( .A(\mem<10><4> ), .B(n984), .Y(n265) );
  OAI21X1 U480 ( .A(n1041), .B(n983), .C(n266), .Y(n788) );
  NAND2X1 U481 ( .A(\mem<10><5> ), .B(n984), .Y(n266) );
  OAI21X1 U482 ( .A(n1042), .B(n983), .C(n267), .Y(n789) );
  NAND2X1 U483 ( .A(\mem<10><6> ), .B(n984), .Y(n267) );
  OAI21X1 U484 ( .A(n1043), .B(n983), .C(n268), .Y(n790) );
  NAND2X1 U485 ( .A(\mem<10><7> ), .B(n984), .Y(n268) );
  NAND3X1 U486 ( .A(n111), .B(n48), .C(n228), .Y(n260) );
  OAI21X1 U487 ( .A(n1028), .B(n982), .C(n270), .Y(n791) );
  NAND2X1 U488 ( .A(\mem<9><0> ), .B(n982), .Y(n270) );
  OAI21X1 U489 ( .A(n1029), .B(n982), .C(n271), .Y(n792) );
  NAND2X1 U490 ( .A(\mem<9><1> ), .B(n982), .Y(n271) );
  OAI21X1 U491 ( .A(n1030), .B(n982), .C(n272), .Y(n793) );
  NAND2X1 U492 ( .A(\mem<9><2> ), .B(n982), .Y(n272) );
  OAI21X1 U493 ( .A(n1031), .B(n982), .C(n273), .Y(n794) );
  NAND2X1 U494 ( .A(\mem<9><3> ), .B(n982), .Y(n273) );
  OAI21X1 U495 ( .A(n1032), .B(n982), .C(n274), .Y(n795) );
  NAND2X1 U496 ( .A(\mem<9><4> ), .B(n982), .Y(n274) );
  OAI21X1 U497 ( .A(n1033), .B(n982), .C(n275), .Y(n796) );
  NAND2X1 U498 ( .A(\mem<9><5> ), .B(n982), .Y(n275) );
  OAI21X1 U499 ( .A(n1034), .B(n982), .C(n276), .Y(n797) );
  NAND2X1 U500 ( .A(\mem<9><6> ), .B(n982), .Y(n276) );
  OAI21X1 U501 ( .A(n1035), .B(n982), .C(n277), .Y(n798) );
  NAND2X1 U502 ( .A(\mem<9><7> ), .B(n982), .Y(n277) );
  NAND3X1 U503 ( .A(n973), .B(n48), .C(n278), .Y(n269) );
  OAI21X1 U504 ( .A(n1036), .B(n981), .C(n280), .Y(n799) );
  NAND2X1 U505 ( .A(\mem<8><0> ), .B(n981), .Y(n280) );
  OAI21X1 U506 ( .A(n1037), .B(n980), .C(n281), .Y(n800) );
  NAND2X1 U507 ( .A(\mem<8><1> ), .B(n981), .Y(n281) );
  OAI21X1 U508 ( .A(n1038), .B(n980), .C(n282), .Y(n801) );
  NAND2X1 U509 ( .A(\mem<8><2> ), .B(n981), .Y(n282) );
  OAI21X1 U510 ( .A(n1039), .B(n980), .C(n283), .Y(n802) );
  NAND2X1 U511 ( .A(\mem<8><3> ), .B(n981), .Y(n283) );
  OAI21X1 U512 ( .A(n1040), .B(n980), .C(n284), .Y(n803) );
  NAND2X1 U513 ( .A(\mem<8><4> ), .B(n981), .Y(n284) );
  OAI21X1 U514 ( .A(n1041), .B(n980), .C(n285), .Y(n804) );
  NAND2X1 U515 ( .A(\mem<8><5> ), .B(n981), .Y(n285) );
  OAI21X1 U516 ( .A(n1042), .B(n980), .C(n286), .Y(n805) );
  NAND2X1 U517 ( .A(\mem<8><6> ), .B(n981), .Y(n286) );
  OAI21X1 U518 ( .A(n1043), .B(n980), .C(n287), .Y(n806) );
  NAND2X1 U519 ( .A(\mem<8><7> ), .B(n981), .Y(n287) );
  NAND3X1 U520 ( .A(n111), .B(n48), .C(n248), .Y(n279) );
  OAI21X1 U521 ( .A(n1028), .B(n979), .C(n291), .Y(n807) );
  NAND2X1 U522 ( .A(\mem<7><0> ), .B(n979), .Y(n291) );
  OAI21X1 U523 ( .A(n1029), .B(n979), .C(n292), .Y(n808) );
  NAND2X1 U524 ( .A(\mem<7><1> ), .B(n979), .Y(n292) );
  OAI21X1 U525 ( .A(n1030), .B(n979), .C(n293), .Y(n809) );
  NAND2X1 U526 ( .A(\mem<7><2> ), .B(n979), .Y(n293) );
  OAI21X1 U527 ( .A(n1031), .B(n979), .C(n294), .Y(n810) );
  NAND2X1 U528 ( .A(\mem<7><3> ), .B(n979), .Y(n294) );
  OAI21X1 U529 ( .A(n1032), .B(n979), .C(n295), .Y(n811) );
  NAND2X1 U530 ( .A(\mem<7><4> ), .B(n979), .Y(n295) );
  OAI21X1 U531 ( .A(n1033), .B(n979), .C(n296), .Y(n812) );
  NAND2X1 U532 ( .A(\mem<7><5> ), .B(n979), .Y(n296) );
  OAI21X1 U533 ( .A(n1034), .B(n979), .C(n297), .Y(n813) );
  NAND2X1 U534 ( .A(\mem<7><6> ), .B(n979), .Y(n297) );
  OAI21X1 U535 ( .A(n1035), .B(n979), .C(n298), .Y(n814) );
  NAND2X1 U536 ( .A(\mem<7><7> ), .B(n979), .Y(n298) );
  NAND3X1 U537 ( .A(n973), .B(n48), .C(n299), .Y(n290) );
  OAI21X1 U538 ( .A(n1036), .B(n978), .C(n301), .Y(n815) );
  NAND2X1 U539 ( .A(\mem<6><0> ), .B(n978), .Y(n301) );
  OAI21X1 U540 ( .A(n1037), .B(n978), .C(n302), .Y(n816) );
  NAND2X1 U541 ( .A(\mem<6><1> ), .B(n978), .Y(n302) );
  OAI21X1 U542 ( .A(n1038), .B(n978), .C(n303), .Y(n817) );
  NAND2X1 U543 ( .A(\mem<6><2> ), .B(n978), .Y(n303) );
  OAI21X1 U544 ( .A(n1039), .B(n978), .C(n304), .Y(n818) );
  NAND2X1 U545 ( .A(\mem<6><3> ), .B(n978), .Y(n304) );
  OAI21X1 U546 ( .A(n1040), .B(n978), .C(n305), .Y(n819) );
  NAND2X1 U547 ( .A(\mem<6><4> ), .B(n978), .Y(n305) );
  OAI21X1 U548 ( .A(n1041), .B(n978), .C(n306), .Y(n820) );
  NAND2X1 U549 ( .A(\mem<6><5> ), .B(n978), .Y(n306) );
  OAI21X1 U550 ( .A(n1042), .B(n978), .C(n307), .Y(n821) );
  NAND2X1 U551 ( .A(\mem<6><6> ), .B(n978), .Y(n307) );
  OAI21X1 U552 ( .A(n1043), .B(n978), .C(n308), .Y(n822) );
  NAND2X1 U553 ( .A(\mem<6><7> ), .B(n978), .Y(n308) );
  NAND3X1 U554 ( .A(n969), .B(n48), .C(n228), .Y(n300) );
  OAI21X1 U555 ( .A(n1028), .B(n977), .C(n310), .Y(n823) );
  NAND2X1 U556 ( .A(\mem<5><0> ), .B(n977), .Y(n310) );
  OAI21X1 U557 ( .A(n1029), .B(n977), .C(n311), .Y(n824) );
  NAND2X1 U558 ( .A(\mem<5><1> ), .B(n977), .Y(n311) );
  OAI21X1 U559 ( .A(n1030), .B(n977), .C(n312), .Y(n825) );
  NAND2X1 U560 ( .A(\mem<5><2> ), .B(n977), .Y(n312) );
  OAI21X1 U561 ( .A(n1031), .B(n977), .C(n313), .Y(n826) );
  NAND2X1 U562 ( .A(\mem<5><3> ), .B(n977), .Y(n313) );
  OAI21X1 U563 ( .A(n1032), .B(n977), .C(n314), .Y(n827) );
  NAND2X1 U564 ( .A(\mem<5><4> ), .B(n977), .Y(n314) );
  OAI21X1 U565 ( .A(n1033), .B(n977), .C(n315), .Y(n828) );
  NAND2X1 U566 ( .A(\mem<5><5> ), .B(n977), .Y(n315) );
  OAI21X1 U567 ( .A(n1034), .B(n977), .C(n316), .Y(n829) );
  NAND2X1 U568 ( .A(\mem<5><6> ), .B(n977), .Y(n316) );
  OAI21X1 U569 ( .A(n1035), .B(n977), .C(n317), .Y(n830) );
  NAND2X1 U570 ( .A(\mem<5><7> ), .B(n977), .Y(n317) );
  NAND3X1 U571 ( .A(n973), .B(n48), .C(n318), .Y(n309) );
  OAI21X1 U572 ( .A(n1036), .B(n976), .C(n320), .Y(n831) );
  NAND2X1 U573 ( .A(\mem<4><0> ), .B(n976), .Y(n320) );
  OAI21X1 U574 ( .A(n1037), .B(n976), .C(n321), .Y(n832) );
  NAND2X1 U575 ( .A(\mem<4><1> ), .B(n976), .Y(n321) );
  OAI21X1 U576 ( .A(n1038), .B(n976), .C(n322), .Y(n833) );
  NAND2X1 U577 ( .A(\mem<4><2> ), .B(n976), .Y(n322) );
  OAI21X1 U578 ( .A(n1039), .B(n976), .C(n323), .Y(n834) );
  NAND2X1 U579 ( .A(\mem<4><3> ), .B(n976), .Y(n323) );
  OAI21X1 U580 ( .A(n1040), .B(n976), .C(n324), .Y(n835) );
  NAND2X1 U581 ( .A(\mem<4><4> ), .B(n976), .Y(n324) );
  OAI21X1 U582 ( .A(n1041), .B(n976), .C(n325), .Y(n836) );
  NAND2X1 U583 ( .A(\mem<4><5> ), .B(n976), .Y(n325) );
  OAI21X1 U584 ( .A(n1042), .B(n976), .C(n326), .Y(n837) );
  NAND2X1 U585 ( .A(\mem<4><6> ), .B(n976), .Y(n326) );
  OAI21X1 U586 ( .A(n1043), .B(n976), .C(n327), .Y(n838) );
  NAND2X1 U587 ( .A(\mem<4><7> ), .B(n976), .Y(n327) );
  NAND3X1 U588 ( .A(n969), .B(n48), .C(n248), .Y(n319) );
  OAI21X1 U590 ( .A(n1028), .B(n975), .C(n330), .Y(n839) );
  NAND2X1 U591 ( .A(\mem<3><0> ), .B(n975), .Y(n330) );
  OAI21X1 U592 ( .A(n1029), .B(n975), .C(n331), .Y(n840) );
  NAND2X1 U593 ( .A(\mem<3><1> ), .B(n975), .Y(n331) );
  OAI21X1 U594 ( .A(n1030), .B(n975), .C(n332), .Y(n841) );
  NAND2X1 U595 ( .A(\mem<3><2> ), .B(n975), .Y(n332) );
  OAI21X1 U596 ( .A(n1031), .B(n975), .C(n333), .Y(n842) );
  NAND2X1 U597 ( .A(\mem<3><3> ), .B(n975), .Y(n333) );
  OAI21X1 U598 ( .A(n1032), .B(n975), .C(n334), .Y(n843) );
  NAND2X1 U599 ( .A(\mem<3><4> ), .B(n975), .Y(n334) );
  OAI21X1 U600 ( .A(n1033), .B(n975), .C(n335), .Y(n844) );
  NAND2X1 U601 ( .A(\mem<3><5> ), .B(n975), .Y(n335) );
  OAI21X1 U602 ( .A(n1034), .B(n975), .C(n336), .Y(n845) );
  NAND2X1 U603 ( .A(\mem<3><6> ), .B(n975), .Y(n336) );
  OAI21X1 U604 ( .A(n1035), .B(n975), .C(n337), .Y(n846) );
  NAND2X1 U605 ( .A(\mem<3><7> ), .B(n975), .Y(n337) );
  NAND3X1 U606 ( .A(n973), .B(n48), .C(n338), .Y(n329) );
  OAI21X1 U607 ( .A(n1036), .B(n974), .C(n340), .Y(n847) );
  NAND2X1 U608 ( .A(\mem<2><0> ), .B(n974), .Y(n340) );
  OAI21X1 U609 ( .A(n1037), .B(n974), .C(n341), .Y(n848) );
  NAND2X1 U610 ( .A(\mem<2><1> ), .B(n974), .Y(n341) );
  OAI21X1 U611 ( .A(n1038), .B(n974), .C(n342), .Y(n849) );
  NAND2X1 U612 ( .A(\mem<2><2> ), .B(n974), .Y(n342) );
  OAI21X1 U613 ( .A(n1039), .B(n974), .C(n343), .Y(n850) );
  NAND2X1 U614 ( .A(\mem<2><3> ), .B(n974), .Y(n343) );
  OAI21X1 U615 ( .A(n1040), .B(n974), .C(n344), .Y(n851) );
  NAND2X1 U616 ( .A(\mem<2><4> ), .B(n974), .Y(n344) );
  OAI21X1 U617 ( .A(n1041), .B(n974), .C(n345), .Y(n852) );
  NAND2X1 U618 ( .A(\mem<2><5> ), .B(n974), .Y(n345) );
  OAI21X1 U619 ( .A(n1042), .B(n974), .C(n346), .Y(n853) );
  NAND2X1 U620 ( .A(\mem<2><6> ), .B(n974), .Y(n346) );
  OAI21X1 U621 ( .A(n1043), .B(n974), .C(n347), .Y(n854) );
  NAND2X1 U622 ( .A(\mem<2><7> ), .B(n974), .Y(n347) );
  NAND3X1 U623 ( .A(n967), .B(n48), .C(n228), .Y(n339) );
  OAI21X1 U624 ( .A(n1028), .B(n8), .C(n349), .Y(n855) );
  NAND2X1 U625 ( .A(\mem<1><0> ), .B(n8), .Y(n349) );
  OAI21X1 U626 ( .A(n1029), .B(n8), .C(n350), .Y(n856) );
  NAND2X1 U627 ( .A(\mem<1><1> ), .B(n8), .Y(n350) );
  OAI21X1 U628 ( .A(n1030), .B(n8), .C(n351), .Y(n857) );
  NAND2X1 U629 ( .A(\mem<1><2> ), .B(n8), .Y(n351) );
  OAI21X1 U630 ( .A(n1031), .B(n8), .C(n352), .Y(n858) );
  NAND2X1 U631 ( .A(\mem<1><3> ), .B(n8), .Y(n352) );
  OAI21X1 U632 ( .A(n1032), .B(n8), .C(n353), .Y(n859) );
  NAND2X1 U633 ( .A(\mem<1><4> ), .B(n8), .Y(n353) );
  OAI21X1 U634 ( .A(n1033), .B(n8), .C(n354), .Y(n860) );
  NAND2X1 U635 ( .A(\mem<1><5> ), .B(n8), .Y(n354) );
  OAI21X1 U636 ( .A(n1034), .B(n8), .C(n355), .Y(n861) );
  NAND2X1 U637 ( .A(\mem<1><6> ), .B(n8), .Y(n355) );
  OAI21X1 U638 ( .A(n1035), .B(n8), .C(n356), .Y(n862) );
  NAND2X1 U639 ( .A(\mem<1><7> ), .B(n8), .Y(n356) );
  NOR2X1 U641 ( .A(n965), .B(\addr_1c<4> ), .Y(n59) );
  OAI21X1 U642 ( .A(n1036), .B(n972), .C(n359), .Y(n863) );
  NAND2X1 U643 ( .A(\mem<0><0> ), .B(n972), .Y(n359) );
  OAI21X1 U644 ( .A(n1037), .B(n972), .C(n360), .Y(n864) );
  NAND2X1 U645 ( .A(\mem<0><1> ), .B(n972), .Y(n360) );
  OAI21X1 U646 ( .A(n1038), .B(n972), .C(n361), .Y(n865) );
  NAND2X1 U647 ( .A(\mem<0><2> ), .B(n972), .Y(n361) );
  OAI21X1 U648 ( .A(n1039), .B(n972), .C(n362), .Y(n866) );
  NAND2X1 U649 ( .A(\mem<0><3> ), .B(n972), .Y(n362) );
  OAI21X1 U650 ( .A(n1040), .B(n972), .C(n363), .Y(n867) );
  NAND2X1 U651 ( .A(\mem<0><4> ), .B(n972), .Y(n363) );
  OAI21X1 U652 ( .A(n1041), .B(n972), .C(n364), .Y(n868) );
  NAND2X1 U653 ( .A(\mem<0><5> ), .B(n972), .Y(n364) );
  OAI21X1 U654 ( .A(n1042), .B(n972), .C(n365), .Y(n869) );
  NAND2X1 U655 ( .A(\mem<0><6> ), .B(n972), .Y(n365) );
  OAI21X1 U656 ( .A(n1043), .B(n972), .C(n366), .Y(n870) );
  NAND2X1 U657 ( .A(\mem<0><7> ), .B(n972), .Y(n366) );
  NAND3X1 U658 ( .A(n967), .B(n48), .C(n248), .Y(n358) );
  NOR3X1 U661 ( .A(n370), .B(\addr_1c<7> ), .C(\addr_1c<6> ), .Y(n369) );
  NOR3X1 U662 ( .A(n371), .B(\addr_1c<11> ), .C(\addr_1c<10> ), .Y(n368) );
  AOI21X1 U663 ( .A(n473), .B(n373), .C(n963), .Y(n1046) );
  OAI21X1 U665 ( .A(rd), .B(n374), .C(wr), .Y(n373) );
  NAND3X1 U667 ( .A(n375), .B(n1023), .C(n376), .Y(n374) );
  NOR3X1 U668 ( .A(rd1), .B(rd3), .C(rd2), .Y(n376) );
  NOR2X1 U669 ( .A(wr3), .B(wr2), .Y(n375) );
  AOI21X1 U670 ( .A(n460), .B(n378), .C(n1014), .Y(\data_out_1c<9> ) );
  NOR3X1 U671 ( .A(n2), .B(n380), .C(n4), .Y(n378) );
  AOI22X1 U673 ( .A(\mem<16><1> ), .B(n91), .C(\mem<0><1> ), .D(n248), .Y(n383) );
  AOI22X1 U674 ( .A(\mem<18><1> ), .B(n71), .C(\mem<2><1> ), .D(n228), .Y(n382) );
  AOI22X1 U676 ( .A(\mem<20><1> ), .B(n91), .C(\mem<4><1> ), .D(n248), .Y(n385) );
  AOI22X1 U677 ( .A(\mem<22><1> ), .B(n71), .C(\mem<6><1> ), .D(n228), .Y(n384) );
  AOI22X1 U678 ( .A(n288), .B(n893), .C(n249), .D(n933), .Y(n377) );
  AOI22X1 U680 ( .A(\mem<28><1> ), .B(n91), .C(\mem<12><1> ), .D(n248), .Y(
        n389) );
  AOI22X1 U681 ( .A(\mem<30><1> ), .B(n71), .C(\mem<14><1> ), .D(n228), .Y(
        n388) );
  AOI22X1 U683 ( .A(\mem<24><1> ), .B(n91), .C(\mem<8><1> ), .D(n248), .Y(n391) );
  AOI22X1 U684 ( .A(\mem<26><1> ), .B(n71), .C(\mem<10><1> ), .D(n228), .Y(
        n390) );
  AOI21X1 U685 ( .A(n448), .B(n393), .C(n1014), .Y(\data_out_1c<8> ) );
  NOR3X1 U686 ( .A(n940), .B(n395), .C(n950), .Y(n393) );
  AOI21X1 U687 ( .A(n397), .B(n398), .C(n971), .Y(n396) );
  AOI22X1 U688 ( .A(\mem<16><0> ), .B(n91), .C(\mem<0><0> ), .D(n248), .Y(n398) );
  AOI22X1 U689 ( .A(\mem<18><0> ), .B(n71), .C(\mem<2><0> ), .D(n228), .Y(n397) );
  AOI21X1 U690 ( .A(n399), .B(n400), .C(n970), .Y(n394) );
  AOI22X1 U691 ( .A(\mem<20><0> ), .B(n91), .C(\mem<4><0> ), .D(n248), .Y(n400) );
  AOI22X1 U692 ( .A(\mem<22><0> ), .B(n71), .C(\mem<6><0> ), .D(n228), .Y(n399) );
  AOI22X1 U693 ( .A(n288), .B(n891), .C(n249), .D(n931), .Y(n392) );
  AOI22X1 U695 ( .A(\mem<28><0> ), .B(n91), .C(\mem<12><0> ), .D(n248), .Y(
        n404) );
  AOI22X1 U696 ( .A(\mem<30><0> ), .B(n71), .C(\mem<14><0> ), .D(n228), .Y(
        n403) );
  AOI22X1 U698 ( .A(\mem<24><0> ), .B(n91), .C(\mem<8><0> ), .D(n248), .Y(n406) );
  AOI22X1 U699 ( .A(\mem<26><0> ), .B(n71), .C(\mem<10><0> ), .D(n228), .Y(
        n405) );
  OAI21X1 U700 ( .A(n23), .B(n50), .C(rd1), .Y(n407) );
  AOI22X1 U702 ( .A(\mem<17><7> ), .B(n199), .C(\mem<19><7> ), .D(n179), .Y(
        n414) );
  AOI22X1 U703 ( .A(\mem<21><7> ), .B(n160), .C(\mem<23><7> ), .D(n140), .Y(
        n413) );
  AOI22X1 U704 ( .A(\mem<25><7> ), .B(n121), .C(\mem<27><7> ), .D(n101), .Y(
        n411) );
  AOI22X1 U705 ( .A(\mem<29><7> ), .B(n81), .C(\mem<31><7> ), .D(n60), .Y(n410) );
  AOI22X1 U707 ( .A(\mem<1><7> ), .B(n357), .C(\mem<3><7> ), .D(n338), .Y(n419) );
  AOI22X1 U708 ( .A(\mem<5><7> ), .B(n318), .C(\mem<7><7> ), .D(n299), .Y(n418) );
  AOI22X1 U709 ( .A(\mem<9><7> ), .B(n278), .C(\mem<11><7> ), .D(n259), .Y(
        n416) );
  AOI22X1 U710 ( .A(\mem<13><7> ), .B(n238), .C(\mem<15><7> ), .D(n218), .Y(
        n415) );
  OAI21X1 U711 ( .A(n21), .B(n37), .C(rd1), .Y(n420) );
  AOI22X1 U713 ( .A(\mem<17><6> ), .B(n199), .C(\mem<19><6> ), .D(n179), .Y(
        n427) );
  AOI22X1 U714 ( .A(\mem<21><6> ), .B(n160), .C(\mem<23><6> ), .D(n140), .Y(
        n426) );
  AOI22X1 U715 ( .A(\mem<25><6> ), .B(n121), .C(\mem<27><6> ), .D(n101), .Y(
        n424) );
  AOI22X1 U716 ( .A(\mem<29><6> ), .B(n81), .C(\mem<31><6> ), .D(n60), .Y(n423) );
  AOI22X1 U718 ( .A(\mem<1><6> ), .B(n357), .C(\mem<3><6> ), .D(n338), .Y(n432) );
  AOI22X1 U719 ( .A(\mem<5><6> ), .B(n318), .C(\mem<7><6> ), .D(n299), .Y(n431) );
  AOI22X1 U720 ( .A(\mem<9><6> ), .B(n278), .C(\mem<11><6> ), .D(n259), .Y(
        n429) );
  AOI22X1 U721 ( .A(\mem<13><6> ), .B(n238), .C(\mem<15><6> ), .D(n218), .Y(
        n428) );
  OAI21X1 U722 ( .A(n19), .B(n35), .C(rd1), .Y(n433) );
  AOI22X1 U724 ( .A(\mem<17><5> ), .B(n199), .C(\mem<19><5> ), .D(n179), .Y(
        n440) );
  AOI22X1 U725 ( .A(\mem<21><5> ), .B(n160), .C(\mem<23><5> ), .D(n140), .Y(
        n439) );
  AOI22X1 U726 ( .A(\mem<25><5> ), .B(n121), .C(\mem<27><5> ), .D(n101), .Y(
        n437) );
  AOI22X1 U727 ( .A(\mem<29><5> ), .B(n81), .C(\mem<31><5> ), .D(n60), .Y(n436) );
  AOI22X1 U729 ( .A(\mem<1><5> ), .B(n357), .C(\mem<3><5> ), .D(n338), .Y(n445) );
  AOI22X1 U730 ( .A(\mem<5><5> ), .B(n318), .C(\mem<7><5> ), .D(n299), .Y(n444) );
  AOI22X1 U731 ( .A(\mem<9><5> ), .B(n278), .C(\mem<11><5> ), .D(n259), .Y(
        n442) );
  AOI22X1 U732 ( .A(\mem<13><5> ), .B(n238), .C(\mem<15><5> ), .D(n218), .Y(
        n441) );
  OAI21X1 U733 ( .A(n17), .B(n33), .C(rd1), .Y(n446) );
  AOI22X1 U735 ( .A(\mem<17><4> ), .B(n199), .C(\mem<19><4> ), .D(n179), .Y(
        n453) );
  AOI22X1 U736 ( .A(\mem<21><4> ), .B(n160), .C(\mem<23><4> ), .D(n140), .Y(
        n452) );
  AOI22X1 U737 ( .A(\mem<25><4> ), .B(n121), .C(\mem<27><4> ), .D(n101), .Y(
        n450) );
  AOI22X1 U738 ( .A(\mem<29><4> ), .B(n81), .C(\mem<31><4> ), .D(n60), .Y(n449) );
  AOI22X1 U740 ( .A(\mem<1><4> ), .B(n357), .C(\mem<3><4> ), .D(n338), .Y(n458) );
  AOI22X1 U741 ( .A(\mem<5><4> ), .B(n318), .C(\mem<7><4> ), .D(n299), .Y(n457) );
  AOI22X1 U742 ( .A(\mem<9><4> ), .B(n278), .C(\mem<11><4> ), .D(n259), .Y(
        n455) );
  AOI22X1 U743 ( .A(\mem<13><4> ), .B(n238), .C(\mem<15><4> ), .D(n218), .Y(
        n454) );
  OAI21X1 U744 ( .A(n15), .B(n31), .C(rd1), .Y(n459) );
  AOI22X1 U746 ( .A(\mem<17><3> ), .B(n199), .C(\mem<19><3> ), .D(n179), .Y(
        n466) );
  AOI22X1 U747 ( .A(\mem<21><3> ), .B(n160), .C(\mem<23><3> ), .D(n140), .Y(
        n465) );
  AOI22X1 U748 ( .A(\mem<25><3> ), .B(n121), .C(\mem<27><3> ), .D(n101), .Y(
        n463) );
  AOI22X1 U749 ( .A(\mem<29><3> ), .B(n81), .C(\mem<31><3> ), .D(n60), .Y(n462) );
  AOI22X1 U751 ( .A(\mem<1><3> ), .B(n357), .C(\mem<3><3> ), .D(n338), .Y(n471) );
  AOI22X1 U752 ( .A(\mem<5><3> ), .B(n318), .C(\mem<7><3> ), .D(n299), .Y(n470) );
  AOI22X1 U753 ( .A(\mem<9><3> ), .B(n278), .C(\mem<11><3> ), .D(n259), .Y(
        n468) );
  AOI22X1 U754 ( .A(\mem<13><3> ), .B(n238), .C(\mem<15><3> ), .D(n218), .Y(
        n467) );
  OAI21X1 U755 ( .A(n13), .B(n29), .C(rd1), .Y(n472) );
  AOI22X1 U757 ( .A(\mem<17><2> ), .B(n199), .C(\mem<19><2> ), .D(n179), .Y(
        n479) );
  AOI22X1 U758 ( .A(\mem<21><2> ), .B(n160), .C(\mem<23><2> ), .D(n140), .Y(
        n478) );
  AOI22X1 U759 ( .A(\mem<25><2> ), .B(n121), .C(\mem<27><2> ), .D(n101), .Y(
        n476) );
  AOI22X1 U760 ( .A(\mem<29><2> ), .B(n81), .C(\mem<31><2> ), .D(n60), .Y(n475) );
  AOI22X1 U762 ( .A(\mem<1><2> ), .B(n357), .C(\mem<3><2> ), .D(n338), .Y(n484) );
  AOI22X1 U763 ( .A(\mem<5><2> ), .B(n318), .C(\mem<7><2> ), .D(n299), .Y(n483) );
  AOI22X1 U764 ( .A(\mem<9><2> ), .B(n278), .C(\mem<11><2> ), .D(n259), .Y(
        n481) );
  AOI22X1 U765 ( .A(\mem<13><2> ), .B(n238), .C(\mem<15><2> ), .D(n218), .Y(
        n480) );
  OAI21X1 U766 ( .A(n11), .B(n27), .C(rd1), .Y(n485) );
  AOI22X1 U768 ( .A(\mem<17><1> ), .B(n199), .C(\mem<19><1> ), .D(n179), .Y(
        n492) );
  AOI22X1 U769 ( .A(\mem<21><1> ), .B(n160), .C(\mem<23><1> ), .D(n140), .Y(
        n491) );
  AOI22X1 U770 ( .A(\mem<25><1> ), .B(n121), .C(\mem<27><1> ), .D(n101), .Y(
        n489) );
  AOI22X1 U771 ( .A(\mem<29><1> ), .B(n81), .C(\mem<31><1> ), .D(n60), .Y(n488) );
  AOI22X1 U773 ( .A(\mem<1><1> ), .B(n357), .C(\mem<3><1> ), .D(n338), .Y(n497) );
  AOI22X1 U774 ( .A(\mem<5><1> ), .B(n318), .C(\mem<7><1> ), .D(n299), .Y(n496) );
  AOI22X1 U775 ( .A(\mem<9><1> ), .B(n278), .C(\mem<11><1> ), .D(n259), .Y(
        n494) );
  AOI22X1 U776 ( .A(\mem<13><1> ), .B(n238), .C(\mem<15><1> ), .D(n218), .Y(
        n493) );
  AOI21X1 U777 ( .A(n447), .B(n499), .C(n1014), .Y(\data_out_1c<15> ) );
  NOR3X1 U778 ( .A(n939), .B(n501), .C(n949), .Y(n499) );
  AOI21X1 U779 ( .A(n503), .B(n504), .C(n971), .Y(n502) );
  AOI22X1 U780 ( .A(\mem<16><7> ), .B(n91), .C(\mem<0><7> ), .D(n248), .Y(n504) );
  AOI22X1 U781 ( .A(\mem<18><7> ), .B(n71), .C(\mem<2><7> ), .D(n228), .Y(n503) );
  AOI21X1 U782 ( .A(n505), .B(n506), .C(n970), .Y(n500) );
  AOI22X1 U783 ( .A(\mem<20><7> ), .B(n91), .C(\mem<4><7> ), .D(n248), .Y(n506) );
  AOI22X1 U784 ( .A(\mem<22><7> ), .B(n71), .C(\mem<6><7> ), .D(n228), .Y(n505) );
  AOI22X1 U785 ( .A(n288), .B(n889), .C(n249), .D(n929), .Y(n498) );
  AOI22X1 U787 ( .A(\mem<28><7> ), .B(n91), .C(\mem<12><7> ), .D(n248), .Y(
        n510) );
  AOI22X1 U788 ( .A(\mem<30><7> ), .B(n71), .C(\mem<14><7> ), .D(n228), .Y(
        n509) );
  AOI22X1 U790 ( .A(\mem<24><7> ), .B(n91), .C(\mem<8><7> ), .D(n248), .Y(n512) );
  AOI22X1 U791 ( .A(\mem<26><7> ), .B(n71), .C(\mem<10><7> ), .D(n228), .Y(
        n511) );
  AOI21X1 U792 ( .A(n435), .B(n514), .C(n1014), .Y(\data_out_1c<14> ) );
  NOR3X1 U793 ( .A(n938), .B(n516), .C(n948), .Y(n514) );
  AOI21X1 U794 ( .A(n518), .B(n519), .C(n971), .Y(n517) );
  AOI22X1 U795 ( .A(\mem<16><6> ), .B(n91), .C(\mem<0><6> ), .D(n248), .Y(n519) );
  AOI22X1 U796 ( .A(\mem<18><6> ), .B(n71), .C(\mem<2><6> ), .D(n228), .Y(n518) );
  AOI21X1 U797 ( .A(n520), .B(n521), .C(n970), .Y(n515) );
  AOI22X1 U798 ( .A(\mem<20><6> ), .B(n91), .C(\mem<4><6> ), .D(n248), .Y(n521) );
  AOI22X1 U799 ( .A(\mem<22><6> ), .B(n71), .C(\mem<6><6> ), .D(n228), .Y(n520) );
  AOI22X1 U800 ( .A(n288), .B(n887), .C(n249), .D(n927), .Y(n513) );
  AOI22X1 U802 ( .A(\mem<28><6> ), .B(n91), .C(\mem<12><6> ), .D(n248), .Y(
        n525) );
  AOI22X1 U803 ( .A(\mem<30><6> ), .B(n71), .C(\mem<14><6> ), .D(n228), .Y(
        n524) );
  AOI22X1 U805 ( .A(\mem<24><6> ), .B(n91), .C(\mem<8><6> ), .D(n248), .Y(n527) );
  AOI22X1 U806 ( .A(\mem<26><6> ), .B(n71), .C(\mem<10><6> ), .D(n228), .Y(
        n526) );
  AOI21X1 U807 ( .A(n434), .B(n529), .C(n1014), .Y(\data_out_1c<13> ) );
  NOR3X1 U808 ( .A(n937), .B(n531), .C(n947), .Y(n529) );
  AOI21X1 U809 ( .A(n533), .B(n534), .C(n971), .Y(n532) );
  AOI22X1 U810 ( .A(\mem<16><5> ), .B(n91), .C(\mem<0><5> ), .D(n248), .Y(n534) );
  AOI22X1 U811 ( .A(\mem<18><5> ), .B(n71), .C(\mem<2><5> ), .D(n228), .Y(n533) );
  AOI21X1 U812 ( .A(n535), .B(n536), .C(n970), .Y(n530) );
  AOI22X1 U813 ( .A(\mem<20><5> ), .B(n91), .C(\mem<4><5> ), .D(n248), .Y(n536) );
  AOI22X1 U814 ( .A(\mem<22><5> ), .B(n71), .C(\mem<6><5> ), .D(n228), .Y(n535) );
  AOI22X1 U815 ( .A(n288), .B(n885), .C(n249), .D(n925), .Y(n528) );
  AOI22X1 U817 ( .A(\mem<28><5> ), .B(n91), .C(\mem<12><5> ), .D(n248), .Y(
        n540) );
  AOI22X1 U818 ( .A(\mem<30><5> ), .B(n71), .C(\mem<14><5> ), .D(n228), .Y(
        n539) );
  AOI22X1 U820 ( .A(\mem<24><5> ), .B(n91), .C(\mem<8><5> ), .D(n248), .Y(n542) );
  AOI22X1 U821 ( .A(\mem<26><5> ), .B(n71), .C(\mem<10><5> ), .D(n228), .Y(
        n541) );
  AOI21X1 U822 ( .A(n422), .B(n544), .C(n1014), .Y(\data_out_1c<12> ) );
  NOR3X1 U823 ( .A(n936), .B(n546), .C(n946), .Y(n544) );
  AOI21X1 U824 ( .A(n548), .B(n549), .C(n971), .Y(n547) );
  AOI22X1 U825 ( .A(\mem<16><4> ), .B(n91), .C(\mem<0><4> ), .D(n248), .Y(n549) );
  AOI22X1 U826 ( .A(\mem<18><4> ), .B(n71), .C(\mem<2><4> ), .D(n228), .Y(n548) );
  AOI21X1 U827 ( .A(n550), .B(n551), .C(n970), .Y(n545) );
  AOI22X1 U828 ( .A(\mem<20><4> ), .B(n91), .C(\mem<4><4> ), .D(n248), .Y(n551) );
  AOI22X1 U829 ( .A(\mem<22><4> ), .B(n71), .C(\mem<6><4> ), .D(n228), .Y(n550) );
  AOI22X1 U830 ( .A(n288), .B(n883), .C(n249), .D(n923), .Y(n543) );
  AOI22X1 U832 ( .A(\mem<28><4> ), .B(n91), .C(\mem<12><4> ), .D(n248), .Y(
        n555) );
  AOI22X1 U833 ( .A(\mem<30><4> ), .B(n71), .C(\mem<14><4> ), .D(n228), .Y(
        n554) );
  AOI22X1 U835 ( .A(\mem<24><4> ), .B(n91), .C(\mem<8><4> ), .D(n248), .Y(n557) );
  AOI22X1 U836 ( .A(\mem<26><4> ), .B(n71), .C(\mem<10><4> ), .D(n228), .Y(
        n556) );
  AOI21X1 U837 ( .A(n421), .B(n559), .C(n1014), .Y(\data_out_1c<11> ) );
  NOR3X1 U838 ( .A(n935), .B(n561), .C(n945), .Y(n559) );
  AOI21X1 U839 ( .A(n563), .B(n564), .C(n971), .Y(n562) );
  AOI22X1 U840 ( .A(\mem<16><3> ), .B(n91), .C(\mem<0><3> ), .D(n248), .Y(n564) );
  AOI22X1 U841 ( .A(\mem<18><3> ), .B(n71), .C(\mem<2><3> ), .D(n228), .Y(n563) );
  AOI21X1 U842 ( .A(n565), .B(n566), .C(n970), .Y(n560) );
  AOI22X1 U843 ( .A(\mem<20><3> ), .B(n91), .C(\mem<4><3> ), .D(n248), .Y(n566) );
  AOI22X1 U844 ( .A(\mem<22><3> ), .B(n71), .C(\mem<6><3> ), .D(n228), .Y(n565) );
  AOI22X1 U845 ( .A(n288), .B(n881), .C(n249), .D(n921), .Y(n558) );
  AOI22X1 U847 ( .A(\mem<28><3> ), .B(n91), .C(\mem<12><3> ), .D(n248), .Y(
        n570) );
  AOI22X1 U848 ( .A(\mem<30><3> ), .B(n71), .C(\mem<14><3> ), .D(n228), .Y(
        n569) );
  AOI22X1 U850 ( .A(\mem<24><3> ), .B(n91), .C(\mem<8><3> ), .D(n248), .Y(n572) );
  AOI22X1 U851 ( .A(\mem<26><3> ), .B(n71), .C(\mem<10><3> ), .D(n228), .Y(
        n571) );
  AOI21X1 U852 ( .A(n409), .B(n574), .C(n1014), .Y(\data_out_1c<10> ) );
  NOR3X1 U853 ( .A(n934), .B(n576), .C(n944), .Y(n574) );
  AOI21X1 U854 ( .A(n578), .B(n579), .C(n971), .Y(n577) );
  AOI22X1 U855 ( .A(\mem<16><2> ), .B(n91), .C(\mem<0><2> ), .D(n248), .Y(n579) );
  AOI22X1 U856 ( .A(\mem<18><2> ), .B(n71), .C(\mem<2><2> ), .D(n228), .Y(n578) );
  AOI21X1 U857 ( .A(n580), .B(n581), .C(n970), .Y(n575) );
  AOI22X1 U858 ( .A(\mem<20><2> ), .B(n91), .C(\mem<4><2> ), .D(n248), .Y(n581) );
  AOI22X1 U859 ( .A(\mem<22><2> ), .B(n71), .C(\mem<6><2> ), .D(n228), .Y(n580) );
  AOI22X1 U860 ( .A(n288), .B(n879), .C(n249), .D(n919), .Y(n573) );
  AOI22X1 U862 ( .A(\mem<28><2> ), .B(n91), .C(\mem<12><2> ), .D(n248), .Y(
        n585) );
  AOI22X1 U863 ( .A(\mem<30><2> ), .B(n71), .C(\mem<14><2> ), .D(n228), .Y(
        n584) );
  AOI22X1 U865 ( .A(\mem<24><2> ), .B(n91), .C(\mem<8><2> ), .D(n248), .Y(n587) );
  AOI22X1 U866 ( .A(\mem<26><2> ), .B(n71), .C(\mem<10><2> ), .D(n228), .Y(
        n586) );
  NOR2X1 U867 ( .A(\addr_1c<3> ), .B(\addr_1c<4> ), .Y(n588) );
  NOR2X1 U868 ( .A(n1027), .B(\addr_1c<4> ), .Y(n589) );
  OAI21X1 U869 ( .A(n9), .B(n25), .C(rd1), .Y(n590) );
  AOI22X1 U871 ( .A(\mem<17><0> ), .B(n199), .C(\mem<19><0> ), .D(n179), .Y(
        n597) );
  AOI22X1 U872 ( .A(\mem<21><0> ), .B(n160), .C(\mem<23><0> ), .D(n140), .Y(
        n596) );
  AOI22X1 U873 ( .A(\mem<25><0> ), .B(n121), .C(\mem<27><0> ), .D(n101), .Y(
        n594) );
  AOI22X1 U874 ( .A(\mem<29><0> ), .B(n81), .C(\mem<31><0> ), .D(n60), .Y(n593) );
  AOI22X1 U876 ( .A(\mem<1><0> ), .B(n357), .C(\mem<3><0> ), .D(n338), .Y(n604) );
  NAND2X1 U877 ( .A(n1025), .B(n1026), .Y(n367) );
  AOI22X1 U878 ( .A(\mem<5><0> ), .B(n318), .C(\mem<7><0> ), .D(n299), .Y(n603) );
  NAND2X1 U879 ( .A(\addr_1c<1> ), .B(n1026), .Y(n328) );
  AOI22X1 U880 ( .A(\mem<9><0> ), .B(n278), .C(\mem<11><0> ), .D(n259), .Y(
        n601) );
  AOI22X1 U881 ( .A(\mem<13><0> ), .B(n238), .C(\mem<15><0> ), .D(n218), .Y(
        n600) );
  dff_207 ff0 ( .q(rd1), .d(rd0), .clk(clk), .rst(n1012) );
  dff_206 ff1 ( .q(wr1), .d(wr0), .clk(clk), .rst(n1012) );
  dff_189 \reg0[0]  ( .q(\addr_1c<0> ), .d(\addr<0> ), .clk(clk), .rst(n1012)
         );
  dff_190 \reg0[1]  ( .q(\addr_1c<1> ), .d(\addr<1> ), .clk(clk), .rst(n1012)
         );
  dff_191 \reg0[2]  ( .q(\addr_1c<2> ), .d(\addr<2> ), .clk(clk), .rst(n1012)
         );
  dff_192 \reg0[3]  ( .q(\addr_1c<3> ), .d(\addr<3> ), .clk(clk), .rst(n1012)
         );
  dff_193 \reg0[4]  ( .q(\addr_1c<4> ), .d(\addr<4> ), .clk(clk), .rst(n1012)
         );
  dff_194 \reg0[5]  ( .q(\addr_1c<5> ), .d(\addr<5> ), .clk(clk), .rst(n1012)
         );
  dff_195 \reg0[6]  ( .q(\addr_1c<6> ), .d(\addr<6> ), .clk(clk), .rst(n1012)
         );
  dff_196 \reg0[7]  ( .q(\addr_1c<7> ), .d(\addr<7> ), .clk(clk), .rst(n1012)
         );
  dff_197 \reg0[8]  ( .q(\addr_1c<8> ), .d(\addr<8> ), .clk(clk), .rst(n1012)
         );
  dff_198 \reg0[9]  ( .q(\addr_1c<9> ), .d(\addr<9> ), .clk(clk), .rst(n1012)
         );
  dff_199 \reg0[10]  ( .q(\addr_1c<10> ), .d(\addr<10> ), .clk(clk), .rst(
        n1012) );
  dff_200 \reg0[11]  ( .q(\addr_1c<11> ), .d(\addr<11> ), .clk(clk), .rst(
        n1012) );
  dff_201 \reg0[12]  ( .q(\addr_1c<12> ), .d(\addr<12> ), .clk(clk), .rst(
        n1012) );
  dff_173 \reg1[0]  ( .q(\data_in_1c<0> ), .d(\data_in<0> ), .clk(clk), .rst(
        n1012) );
  dff_174 \reg1[1]  ( .q(\data_in_1c<1> ), .d(\data_in<1> ), .clk(clk), .rst(
        n1012) );
  dff_175 \reg1[2]  ( .q(\data_in_1c<2> ), .d(\data_in<2> ), .clk(clk), .rst(
        n1012) );
  dff_176 \reg1[3]  ( .q(\data_in_1c<3> ), .d(\data_in<3> ), .clk(clk), .rst(
        n1012) );
  dff_177 \reg1[4]  ( .q(\data_in_1c<4> ), .d(\data_in<4> ), .clk(clk), .rst(
        n1012) );
  dff_178 \reg1[5]  ( .q(\data_in_1c<5> ), .d(\data_in<5> ), .clk(clk), .rst(
        n1012) );
  dff_179 \reg1[6]  ( .q(\data_in_1c<6> ), .d(\data_in<6> ), .clk(clk), .rst(
        n1012) );
  dff_180 \reg1[7]  ( .q(\data_in_1c<7> ), .d(\data_in<7> ), .clk(clk), .rst(
        n1012) );
  dff_181 \reg1[8]  ( .q(\data_in_1c<8> ), .d(\data_in<8> ), .clk(clk), .rst(
        n1012) );
  dff_182 \reg1[9]  ( .q(\data_in_1c<9> ), .d(\data_in<9> ), .clk(clk), .rst(
        n1012) );
  dff_183 \reg1[10]  ( .q(\data_in_1c<10> ), .d(\data_in<10> ), .clk(clk), 
        .rst(n1012) );
  dff_184 \reg1[11]  ( .q(\data_in_1c<11> ), .d(\data_in<11> ), .clk(clk), 
        .rst(n1012) );
  dff_185 \reg1[12]  ( .q(\data_in_1c<12> ), .d(\data_in<12> ), .clk(clk), 
        .rst(n1012) );
  dff_186 \reg1[13]  ( .q(\data_in_1c<13> ), .d(\data_in<13> ), .clk(clk), 
        .rst(n1012) );
  dff_187 \reg1[14]  ( .q(\data_in_1c<14> ), .d(\data_in<14> ), .clk(clk), 
        .rst(n1012) );
  dff_188 \reg1[15]  ( .q(\data_in_1c<15> ), .d(\data_in<15> ), .clk(clk), 
        .rst(n1012) );
  dff_157 \reg2[0]  ( .q(\data_out<0> ), .d(n1022), .clk(clk), .rst(n1012) );
  dff_158 \reg2[1]  ( .q(\data_out<1> ), .d(n1021), .clk(clk), .rst(n1012) );
  dff_159 \reg2[2]  ( .q(\data_out<2> ), .d(n1020), .clk(clk), .rst(n1012) );
  dff_160 \reg2[3]  ( .q(\data_out<3> ), .d(n1019), .clk(clk), .rst(n1012) );
  dff_161 \reg2[4]  ( .q(\data_out<4> ), .d(n1018), .clk(clk), .rst(n1012) );
  dff_162 \reg2[5]  ( .q(\data_out<5> ), .d(n1017), .clk(clk), .rst(n1012) );
  dff_163 \reg2[6]  ( .q(\data_out<6> ), .d(n1016), .clk(clk), .rst(n1012) );
  dff_164 \reg2[7]  ( .q(\data_out<7> ), .d(n1015), .clk(clk), .rst(n1012) );
  dff_165 \reg2[8]  ( .q(\data_out<8> ), .d(\data_out_1c<8> ), .clk(clk), 
        .rst(n1012) );
  dff_166 \reg2[9]  ( .q(\data_out<9> ), .d(\data_out_1c<9> ), .clk(clk), 
        .rst(n1012) );
  dff_167 \reg2[10]  ( .q(\data_out<10> ), .d(\data_out_1c<10> ), .clk(clk), 
        .rst(n1012) );
  dff_168 \reg2[11]  ( .q(\data_out<11> ), .d(\data_out_1c<11> ), .clk(clk), 
        .rst(n1012) );
  dff_169 \reg2[12]  ( .q(\data_out<12> ), .d(\data_out_1c<12> ), .clk(clk), 
        .rst(n1012) );
  dff_170 \reg2[13]  ( .q(\data_out<13> ), .d(\data_out_1c<13> ), .clk(clk), 
        .rst(n1012) );
  dff_171 \reg2[14]  ( .q(\data_out<14> ), .d(\data_out_1c<14> ), .clk(clk), 
        .rst(n1012) );
  dff_172 \reg2[15]  ( .q(\data_out<15> ), .d(\data_out_1c<15> ), .clk(clk), 
        .rst(n1012) );
  dff_205 ff2 ( .q(rd2), .d(rd1), .clk(clk), .rst(n1012) );
  dff_204 ff3 ( .q(wr2), .d(wr1), .clk(clk), .rst(n1012) );
  dff_203 ff4 ( .q(rd3), .d(rd2), .clk(clk), .rst(n1012) );
  dff_202 ff5 ( .q(wr3), .d(wr2), .clk(clk), .rst(n1012) );
  INVX1 U2 ( .A(rd), .Y(n1045) );
  OR2X1 U3 ( .A(\addr_1c<5> ), .B(\addr_1c<12> ), .Y(n371) );
  AND2X1 U4 ( .A(\addr_1c<4> ), .B(n357), .Y(n49) );
  INVX1 U5 ( .A(\addr_1c<3> ), .Y(n1027) );
  INVX1 U6 ( .A(\addr_1c<2> ), .Y(n1026) );
  INVX1 U7 ( .A(wr1), .Y(n1023) );
  INVX1 U8 ( .A(\addr_1c<1> ), .Y(n1025) );
  OR2X1 U23 ( .A(\addr_1c<9> ), .B(\addr_1c<8> ), .Y(n370) );
  AND2X1 U24 ( .A(\addr_1c<3> ), .B(\addr_1c<0> ), .Y(n598) );
  AND2X1 U25 ( .A(\addr_1c<3> ), .B(n1024), .Y(n599) );
  AND2X1 U26 ( .A(n249), .B(n964), .Y(n70) );
  AND2X1 U27 ( .A(n288), .B(n964), .Y(n111) );
  AND2X1 U28 ( .A(\addr_1c<0> ), .B(n1027), .Y(n605) );
  AND2X1 U29 ( .A(n1024), .B(n1027), .Y(n606) );
  INVX1 U35 ( .A(\addr_1c<0> ), .Y(n1024) );
  AND2X1 U36 ( .A(\addr_1c<2> ), .B(n1025), .Y(n288) );
  AND2X1 U37 ( .A(\addr_1c<2> ), .B(\addr_1c<1> ), .Y(n249) );
  AND2X1 U38 ( .A(n599), .B(n249), .Y(n81) );
  AND2X1 U39 ( .A(n288), .B(n598), .Y(n101) );
  AND2X1 U40 ( .A(n288), .B(n599), .Y(n121) );
  AND2X1 U41 ( .A(n941), .B(n598), .Y(n140) );
  AND2X1 U42 ( .A(n941), .B(n599), .Y(n160) );
  AND2X1 U43 ( .A(n598), .B(n951), .Y(n179) );
  AND2X1 U44 ( .A(n599), .B(n951), .Y(n199) );
  AND2X1 U46 ( .A(n605), .B(n249), .Y(n218) );
  AND2X1 U47 ( .A(n249), .B(n606), .Y(n238) );
  AND2X1 U48 ( .A(n605), .B(n288), .Y(n259) );
  AND2X1 U49 ( .A(n288), .B(n606), .Y(n278) );
  AND2X1 U50 ( .A(n605), .B(n941), .Y(n299) );
  AND2X1 U51 ( .A(n941), .B(n606), .Y(n318) );
  OR2X1 U52 ( .A(n970), .B(n965), .Y(n968) );
  AND2X1 U53 ( .A(n605), .B(n951), .Y(n338) );
  OR2X1 U54 ( .A(n965), .B(n971), .Y(n966) );
  AND2X1 U55 ( .A(n49), .B(\mem<32><0> ), .Y(n395) );
  AND2X1 U56 ( .A(n49), .B(\mem<32><1> ), .Y(n380) );
  AND2X1 U57 ( .A(n49), .B(\mem<32><2> ), .Y(n576) );
  AND2X1 U58 ( .A(n49), .B(\mem<32><3> ), .Y(n561) );
  AND2X1 U59 ( .A(n49), .B(\mem<32><4> ), .Y(n546) );
  AND2X1 U60 ( .A(n49), .B(\mem<32><5> ), .Y(n531) );
  AND2X1 U61 ( .A(n49), .B(\mem<32><6> ), .Y(n516) );
  AND2X1 U62 ( .A(n49), .B(\mem<32><7> ), .Y(n501) );
  INVX1 U63 ( .A(rd1), .Y(n1014) );
  BUFX2 U64 ( .A(n961), .Y(n1010) );
  BUFX2 U65 ( .A(n961), .Y(n1009) );
  BUFX2 U66 ( .A(n960), .Y(n1007) );
  BUFX2 U67 ( .A(n960), .Y(n1006) );
  BUFX2 U68 ( .A(n959), .Y(n1004) );
  BUFX2 U69 ( .A(n959), .Y(n1003) );
  BUFX2 U70 ( .A(n958), .Y(n1001) );
  BUFX2 U71 ( .A(n958), .Y(n1000) );
  BUFX2 U72 ( .A(n957), .Y(n990) );
  BUFX2 U73 ( .A(n957), .Y(n989) );
  BUFX2 U74 ( .A(n956), .Y(n987) );
  BUFX2 U75 ( .A(n956), .Y(n986) );
  BUFX2 U76 ( .A(n955), .Y(n984) );
  BUFX2 U77 ( .A(n955), .Y(n983) );
  BUFX2 U78 ( .A(n954), .Y(n981) );
  BUFX2 U79 ( .A(n954), .Y(n980) );
  INVX1 U80 ( .A(\data_in_1c<0> ), .Y(n1028) );
  INVX1 U81 ( .A(\data_in_1c<1> ), .Y(n1029) );
  INVX1 U82 ( .A(\data_in_1c<2> ), .Y(n1030) );
  INVX1 U83 ( .A(\data_in_1c<3> ), .Y(n1031) );
  INVX1 U84 ( .A(\data_in_1c<4> ), .Y(n1032) );
  INVX1 U85 ( .A(\data_in_1c<5> ), .Y(n1033) );
  INVX1 U86 ( .A(\data_in_1c<6> ), .Y(n1034) );
  INVX1 U87 ( .A(\data_in_1c<7> ), .Y(n1035) );
  INVX1 U88 ( .A(\data_in_1c<8> ), .Y(n1036) );
  INVX1 U89 ( .A(\data_in_1c<9> ), .Y(n1037) );
  INVX1 U90 ( .A(\data_in_1c<10> ), .Y(n1038) );
  INVX1 U91 ( .A(\data_in_1c<11> ), .Y(n1039) );
  INVX1 U92 ( .A(\data_in_1c<12> ), .Y(n1040) );
  INVX1 U93 ( .A(\data_in_1c<13> ), .Y(n1041) );
  INVX1 U129 ( .A(\data_in_1c<14> ), .Y(n1042) );
  INVX1 U589 ( .A(\data_in_1c<15> ), .Y(n1043) );
  INVX1 U640 ( .A(wr), .Y(n1044) );
  INVX1 U659 ( .A(n590), .Y(n1022) );
  INVX1 U660 ( .A(n485), .Y(n1021) );
  INVX1 U664 ( .A(n472), .Y(n1020) );
  INVX1 U666 ( .A(n459), .Y(n1019) );
  INVX1 U672 ( .A(n446), .Y(n1018) );
  INVX1 U675 ( .A(n433), .Y(n1017) );
  INVX1 U679 ( .A(n420), .Y(n1016) );
  INVX1 U682 ( .A(n407), .Y(n1015) );
  INVX1 U694 ( .A(rst), .Y(n1013) );
  INVX2 U697 ( .A(n1013), .Y(n1012) );
  AND2X1 U701 ( .A(wr1), .B(n1013), .Y(n48) );
  AND2X1 U706 ( .A(n387), .B(n372), .Y(n1) );
  INVX1 U712 ( .A(n1), .Y(n2) );
  AND2X1 U717 ( .A(n402), .B(n381), .Y(n3) );
  INVX1 U723 ( .A(n3), .Y(n4) );
  AND2X1 U728 ( .A(n60), .B(n189), .Y(n5) );
  INVX1 U734 ( .A(n5), .Y(n6) );
  AND2X1 U739 ( .A(n973), .B(n289), .Y(n7) );
  INVX1 U745 ( .A(n7), .Y(n8) );
  OR2X1 U750 ( .A(n487), .B(n10), .Y(n9) );
  OR2X1 U756 ( .A(n474), .B(n486), .Y(n10) );
  OR2X1 U761 ( .A(n522), .B(n12), .Y(n11) );
  OR2X1 U767 ( .A(n507), .B(n508), .Y(n12) );
  OR2X1 U772 ( .A(n538), .B(n14), .Y(n13) );
  OR2X1 U786 ( .A(n523), .B(n537), .Y(n14) );
  OR2X1 U789 ( .A(n567), .B(n16), .Y(n15) );
  OR2X1 U801 ( .A(n552), .B(n553), .Y(n16) );
  OR2X1 U804 ( .A(n583), .B(n18), .Y(n17) );
  OR2X1 U816 ( .A(n568), .B(n582), .Y(n18) );
  OR2X1 U819 ( .A(n871), .B(n20), .Y(n19) );
  OR2X1 U831 ( .A(n591), .B(n592), .Y(n20) );
  OR2X1 U834 ( .A(n874), .B(n22), .Y(n21) );
  OR2X1 U846 ( .A(n872), .B(n873), .Y(n22) );
  OR2X1 U849 ( .A(n877), .B(n24), .Y(n23) );
  OR2X1 U861 ( .A(n875), .B(n876), .Y(n24) );
  OR2X1 U864 ( .A(n896), .B(n26), .Y(n25) );
  OR2X1 U870 ( .A(n894), .B(n895), .Y(n26) );
  OR2X1 U875 ( .A(n899), .B(n28), .Y(n27) );
  OR2X1 U882 ( .A(n897), .B(n898), .Y(n28) );
  OR2X1 U883 ( .A(n902), .B(n30), .Y(n29) );
  OR2X1 U884 ( .A(n900), .B(n901), .Y(n30) );
  OR2X1 U885 ( .A(n905), .B(n32), .Y(n31) );
  OR2X1 U886 ( .A(n903), .B(n904), .Y(n32) );
  OR2X1 U887 ( .A(n908), .B(n34), .Y(n33) );
  OR2X1 U888 ( .A(n906), .B(n907), .Y(n34) );
  OR2X1 U889 ( .A(n911), .B(n36), .Y(n35) );
  OR2X1 U890 ( .A(n909), .B(n910), .Y(n36) );
  OR2X1 U891 ( .A(n914), .B(n38), .Y(n37) );
  OR2X1 U892 ( .A(n912), .B(n913), .Y(n38) );
  OR2X1 U893 ( .A(n917), .B(n150), .Y(n50) );
  OR2X1 U894 ( .A(n915), .B(n916), .Y(n150) );
  AND2X1 U895 ( .A(n973), .B(n48), .Y(n189) );
  AND2X1 U896 ( .A(n48), .B(n357), .Y(n289) );
  AND2X1 U897 ( .A(n941), .B(n943), .Y(n348) );
  INVX1 U898 ( .A(n348), .Y(n372) );
  AND2X1 U899 ( .A(n951), .B(n953), .Y(n379) );
  INVX1 U900 ( .A(n379), .Y(n381) );
  AND2X1 U901 ( .A(n941), .B(n942), .Y(n386) );
  INVX1 U902 ( .A(n386), .Y(n387) );
  AND2X1 U903 ( .A(n951), .B(n952), .Y(n401) );
  INVX1 U904 ( .A(n401), .Y(n402) );
  BUFX2 U905 ( .A(n1046), .Y(err) );
  BUFX2 U906 ( .A(n573), .Y(n409) );
  BUFX2 U907 ( .A(n558), .Y(n421) );
  BUFX2 U908 ( .A(n543), .Y(n422) );
  BUFX2 U909 ( .A(n528), .Y(n434) );
  BUFX2 U910 ( .A(n513), .Y(n435) );
  BUFX2 U911 ( .A(n498), .Y(n447) );
  BUFX2 U912 ( .A(n392), .Y(n448) );
  BUFX2 U913 ( .A(n377), .Y(n460) );
  AND2X2 U914 ( .A(rd), .B(n374), .Y(n461) );
  INVX1 U915 ( .A(n461), .Y(n473) );
  INVX1 U916 ( .A(n602), .Y(n474) );
  INVX1 U917 ( .A(n601), .Y(n486) );
  INVX1 U918 ( .A(n600), .Y(n487) );
  INVX1 U919 ( .A(n495), .Y(n507) );
  INVX1 U920 ( .A(n494), .Y(n508) );
  INVX1 U921 ( .A(n493), .Y(n522) );
  INVX1 U922 ( .A(n482), .Y(n523) );
  INVX1 U923 ( .A(n481), .Y(n537) );
  INVX1 U924 ( .A(n480), .Y(n538) );
  INVX1 U925 ( .A(n469), .Y(n552) );
  INVX1 U926 ( .A(n468), .Y(n553) );
  INVX1 U927 ( .A(n467), .Y(n567) );
  INVX1 U928 ( .A(n456), .Y(n568) );
  INVX1 U929 ( .A(n455), .Y(n582) );
  INVX1 U930 ( .A(n454), .Y(n583) );
  INVX1 U931 ( .A(n443), .Y(n591) );
  INVX1 U932 ( .A(n442), .Y(n592) );
  INVX1 U933 ( .A(n441), .Y(n871) );
  INVX1 U934 ( .A(n430), .Y(n872) );
  INVX1 U935 ( .A(n429), .Y(n873) );
  INVX1 U936 ( .A(n428), .Y(n874) );
  INVX1 U937 ( .A(n417), .Y(n875) );
  INVX1 U938 ( .A(n416), .Y(n876) );
  INVX1 U939 ( .A(n415), .Y(n877) );
  AND2X2 U940 ( .A(n586), .B(n587), .Y(n878) );
  INVX1 U941 ( .A(n878), .Y(n879) );
  AND2X2 U942 ( .A(n571), .B(n572), .Y(n880) );
  INVX1 U943 ( .A(n880), .Y(n881) );
  AND2X2 U944 ( .A(n556), .B(n557), .Y(n882) );
  INVX1 U945 ( .A(n882), .Y(n883) );
  AND2X2 U946 ( .A(n541), .B(n542), .Y(n884) );
  INVX1 U947 ( .A(n884), .Y(n885) );
  AND2X2 U948 ( .A(n526), .B(n527), .Y(n886) );
  INVX1 U949 ( .A(n886), .Y(n887) );
  AND2X2 U950 ( .A(n511), .B(n512), .Y(n888) );
  INVX1 U951 ( .A(n888), .Y(n889) );
  AND2X2 U952 ( .A(n405), .B(n406), .Y(n890) );
  INVX1 U953 ( .A(n890), .Y(n891) );
  AND2X2 U954 ( .A(n390), .B(n391), .Y(n892) );
  INVX1 U955 ( .A(n892), .Y(n893) );
  INVX1 U956 ( .A(n595), .Y(n894) );
  INVX1 U957 ( .A(n594), .Y(n895) );
  INVX1 U958 ( .A(n593), .Y(n896) );
  INVX1 U959 ( .A(n490), .Y(n897) );
  INVX1 U960 ( .A(n489), .Y(n898) );
  INVX1 U961 ( .A(n488), .Y(n899) );
  INVX1 U962 ( .A(n477), .Y(n900) );
  INVX1 U963 ( .A(n476), .Y(n901) );
  INVX1 U964 ( .A(n475), .Y(n902) );
  INVX1 U965 ( .A(n464), .Y(n903) );
  INVX1 U966 ( .A(n463), .Y(n904) );
  INVX1 U967 ( .A(n462), .Y(n905) );
  INVX1 U968 ( .A(n451), .Y(n906) );
  INVX1 U969 ( .A(n450), .Y(n907) );
  INVX1 U970 ( .A(n449), .Y(n908) );
  INVX1 U971 ( .A(n438), .Y(n909) );
  INVX1 U972 ( .A(n437), .Y(n910) );
  INVX1 U973 ( .A(n436), .Y(n911) );
  INVX1 U974 ( .A(n425), .Y(n912) );
  INVX1 U975 ( .A(n424), .Y(n913) );
  INVX1 U976 ( .A(n423), .Y(n914) );
  INVX1 U977 ( .A(n412), .Y(n915) );
  INVX1 U978 ( .A(n411), .Y(n916) );
  INVX1 U979 ( .A(n410), .Y(n917) );
  AND2X2 U980 ( .A(n584), .B(n585), .Y(n918) );
  INVX1 U981 ( .A(n918), .Y(n919) );
  AND2X2 U982 ( .A(n569), .B(n570), .Y(n920) );
  INVX1 U983 ( .A(n920), .Y(n921) );
  AND2X2 U984 ( .A(n554), .B(n555), .Y(n922) );
  INVX1 U985 ( .A(n922), .Y(n923) );
  AND2X2 U986 ( .A(n539), .B(n540), .Y(n924) );
  INVX1 U987 ( .A(n924), .Y(n925) );
  AND2X2 U988 ( .A(n524), .B(n525), .Y(n926) );
  INVX1 U989 ( .A(n926), .Y(n927) );
  AND2X2 U990 ( .A(n509), .B(n510), .Y(n928) );
  INVX1 U991 ( .A(n928), .Y(n929) );
  AND2X2 U992 ( .A(n403), .B(n404), .Y(n930) );
  INVX1 U993 ( .A(n930), .Y(n931) );
  AND2X2 U994 ( .A(n388), .B(n389), .Y(n932) );
  INVX1 U995 ( .A(n932), .Y(n933) );
  BUFX2 U996 ( .A(n575), .Y(n934) );
  BUFX2 U997 ( .A(n560), .Y(n935) );
  BUFX2 U998 ( .A(n545), .Y(n936) );
  BUFX2 U999 ( .A(n530), .Y(n937) );
  BUFX2 U1000 ( .A(n515), .Y(n938) );
  BUFX2 U1001 ( .A(n500), .Y(n939) );
  BUFX2 U1002 ( .A(n394), .Y(n940) );
  INVX1 U1003 ( .A(n970), .Y(n941) );
  INVX1 U1004 ( .A(n385), .Y(n942) );
  INVX1 U1005 ( .A(n384), .Y(n943) );
  BUFX2 U1006 ( .A(n328), .Y(n970) );
  BUFX2 U1007 ( .A(n577), .Y(n944) );
  BUFX2 U1008 ( .A(n562), .Y(n945) );
  BUFX2 U1009 ( .A(n547), .Y(n946) );
  BUFX2 U1010 ( .A(n532), .Y(n947) );
  BUFX2 U1011 ( .A(n517), .Y(n948) );
  BUFX2 U1012 ( .A(n502), .Y(n949) );
  BUFX2 U1013 ( .A(n396), .Y(n950) );
  INVX1 U1014 ( .A(n971), .Y(n951) );
  INVX1 U1015 ( .A(n383), .Y(n952) );
  INVX1 U1016 ( .A(n382), .Y(n953) );
  BUFX2 U1017 ( .A(n367), .Y(n971) );
  BUFX2 U1018 ( .A(n358), .Y(n972) );
  BUFX2 U1019 ( .A(n339), .Y(n974) );
  BUFX2 U1020 ( .A(n329), .Y(n975) );
  BUFX2 U1021 ( .A(n319), .Y(n976) );
  BUFX2 U1022 ( .A(n309), .Y(n977) );
  BUFX2 U1023 ( .A(n300), .Y(n978) );
  BUFX2 U1024 ( .A(n290), .Y(n979) );
  BUFX2 U1025 ( .A(n269), .Y(n982) );
  BUFX2 U1026 ( .A(n250), .Y(n985) );
  BUFX2 U1027 ( .A(n229), .Y(n988) );
  BUFX2 U1028 ( .A(n209), .Y(n991) );
  BUFX2 U1029 ( .A(n200), .Y(n992) );
  BUFX2 U1030 ( .A(n190), .Y(n993) );
  BUFX2 U1031 ( .A(n180), .Y(n994) );
  BUFX2 U1032 ( .A(n170), .Y(n995) );
  BUFX2 U1033 ( .A(n161), .Y(n996) );
  BUFX2 U1034 ( .A(n151), .Y(n997) );
  BUFX2 U1035 ( .A(n141), .Y(n998) );
  BUFX2 U1036 ( .A(n131), .Y(n999) );
  BUFX2 U1037 ( .A(n112), .Y(n1002) );
  BUFX2 U1038 ( .A(n92), .Y(n1005) );
  BUFX2 U1039 ( .A(n72), .Y(n1008) );
  BUFX2 U1040 ( .A(n59), .Y(n973) );
  AND2X1 U1041 ( .A(n249), .B(n598), .Y(n60) );
  BUFX2 U1042 ( .A(n39), .Y(n1011) );
  BUFX2 U1043 ( .A(n279), .Y(n954) );
  BUFX2 U1044 ( .A(n260), .Y(n955) );
  BUFX2 U1045 ( .A(n239), .Y(n956) );
  BUFX2 U1046 ( .A(n219), .Y(n957) );
  BUFX2 U1047 ( .A(n122), .Y(n958) );
  BUFX2 U1048 ( .A(n102), .Y(n959) );
  BUFX2 U1049 ( .A(n82), .Y(n960) );
  BUFX2 U1050 ( .A(n61), .Y(n961) );
  AND2X1 U1051 ( .A(enable), .B(n1013), .Y(n962) );
  INVX1 U1052 ( .A(n962), .Y(n963) );
  AND2X1 U1053 ( .A(n368), .B(n369), .Y(n964) );
  INVX1 U1054 ( .A(n964), .Y(n965) );
  INVX1 U1055 ( .A(n966), .Y(n967) );
  INVX1 U1056 ( .A(n968), .Y(n969) );
  AND2X1 U1057 ( .A(n951), .B(n606), .Y(n357) );
endmodule


module final_memory_2 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), err, .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<12> , \addr<11> , \addr<10> , \addr<9> , 
        \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , 
        \addr<2> , \addr<1> , \addr<0> }), wr, rd, enable, create_dump, 
    .bank_id({\bank_id<1> , \bank_id<0> }), clk, rst );
  input \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , \addr<12> , \addr<11> ,
         \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> , \addr<5> ,
         \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> , wr, rd, enable,
         create_dump, \bank_id<1> , \bank_id<0> , clk, rst;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , err;
  wire   n1838, rd0, wr0, rd1, wr1, \addr_1c<12> , \addr_1c<11> ,
         \addr_1c<10> , \addr_1c<9> , \addr_1c<8> , \addr_1c<7> , \addr_1c<6> ,
         \addr_1c<5> , \addr_1c<4> , \addr_1c<3> , \addr_1c<2> , \addr_1c<1> ,
         \addr_1c<0> , \data_in_1c<15> , \data_in_1c<14> , \data_in_1c<13> ,
         \data_in_1c<12> , \data_in_1c<11> , \data_in_1c<10> , \data_in_1c<9> ,
         \data_in_1c<8> , \data_in_1c<7> , \data_in_1c<6> , \data_in_1c<5> ,
         \data_in_1c<4> , \data_in_1c<3> , \data_in_1c<2> , \data_in_1c<1> ,
         \data_in_1c<0> , \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> ,
         \mem<0><3> , \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><7> ,
         \mem<1><6> , \mem<1><5> , \mem<1><4> , \mem<1><3> , \mem<1><2> ,
         \mem<1><1> , \mem<1><0> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><7> , \mem<3><6> , \mem<3><5> , \mem<3><4> , \mem<3><3> ,
         \mem<3><2> , \mem<3><1> , \mem<3><0> , \mem<4><7> , \mem<4><6> ,
         \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> , \mem<4><1> ,
         \mem<4><0> , \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> ,
         \mem<5><3> , \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><7> ,
         \mem<6><6> , \mem<6><5> , \mem<6><4> , \mem<6><3> , \mem<6><2> ,
         \mem<6><1> , \mem<6><0> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><7> , \mem<8><6> , \mem<8><5> , \mem<8><4> , \mem<8><3> ,
         \mem<8><2> , \mem<8><1> , \mem<8><0> , \mem<9><7> , \mem<9><6> ,
         \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> , \mem<9><1> ,
         \mem<9><0> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><7> ,
         \mem<11><6> , \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> ,
         \mem<11><1> , \mem<11><0> , \mem<12><7> , \mem<12><6> , \mem<12><5> ,
         \mem<12><4> , \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> ,
         \mem<13><7> , \mem<13><6> , \mem<13><5> , \mem<13><4> , \mem<13><3> ,
         \mem<13><2> , \mem<13><1> , \mem<13><0> , \mem<14><7> , \mem<14><6> ,
         \mem<14><5> , \mem<14><4> , \mem<14><3> , \mem<14><2> , \mem<14><1> ,
         \mem<14><0> , \mem<15><7> , \mem<15><6> , \mem<15><5> , \mem<15><4> ,
         \mem<15><3> , \mem<15><2> , \mem<15><1> , \mem<15><0> , \mem<16><7> ,
         \mem<16><6> , \mem<16><5> , \mem<16><4> , \mem<16><3> , \mem<16><2> ,
         \mem<16><1> , \mem<16><0> , \mem<17><7> , \mem<17><6> , \mem<17><5> ,
         \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> , \mem<17><0> ,
         \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> , \mem<18><3> ,
         \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><7> ,
         \mem<21><6> , \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> ,
         \mem<21><1> , \mem<21><0> , \mem<22><7> , \mem<22><6> , \mem<22><5> ,
         \mem<22><4> , \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> ,
         \mem<23><7> , \mem<23><6> , \mem<23><5> , \mem<23><4> , \mem<23><3> ,
         \mem<23><2> , \mem<23><1> , \mem<23><0> , \mem<24><7> , \mem<24><6> ,
         \mem<24><5> , \mem<24><4> , \mem<24><3> , \mem<24><2> , \mem<24><1> ,
         \mem<24><0> , \mem<25><7> , \mem<25><6> , \mem<25><5> , \mem<25><4> ,
         \mem<25><3> , \mem<25><2> , \mem<25><1> , \mem<25><0> , \mem<26><7> ,
         \mem<26><6> , \mem<26><5> , \mem<26><4> , \mem<26><3> , \mem<26><2> ,
         \mem<26><1> , \mem<26><0> , \mem<27><7> , \mem<27><6> , \mem<27><5> ,
         \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> , \mem<27><0> ,
         \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> , \mem<28><3> ,
         \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><7> ,
         \mem<31><6> , \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> ,
         \mem<31><1> , \mem<31><0> , \mem<32><7> , \mem<32><6> , \mem<32><5> ,
         \mem<32><4> , \mem<32><3> , \mem<32><2> , \mem<32><1> , \mem<32><0> ,
         \data_out_1c<15> , \data_out_1c<14> , \data_out_1c<13> ,
         \data_out_1c<12> , \data_out_1c<11> , \data_out_1c<10> ,
         \data_out_1c<9> , \data_out_1c<8> , rd2, wr2, rd3, wr3, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n50, n150, n189, n289, n348, n372, n379,
         n381, n386, n387, n401, n402, n408, n409, n421, n422, n434, n435,
         n447, n448, n460, n461, n473, n474, n486, n487, n507, n508, n522,
         n523, n537, n538, n552, n553, n567, n568, n582, n583, n591, n592,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837;

  DFFPOSX1 \mem_reg<0><7>  ( .D(n1046), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1047), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1048), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1049), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1050), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1051), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1052), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1053), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1054), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1055), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1056), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1057), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1058), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1059), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1060), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1061), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1062), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1063), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1064), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1065), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1066), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1067), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1068), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1069), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1070), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1071), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1072), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1073), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1074), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1075), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1076), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1077), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1078), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1079), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1080), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1081), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1082), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1083), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1084), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1085), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1086), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1087), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1088), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1089), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1090), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1091), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1092), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1093), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1094), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1095), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1096), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1097), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1098), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1099), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1100), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1101), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1102), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1103), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1104), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1105), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1106), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1107), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1108), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1109), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1110), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1111), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1112), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1113), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1114), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1115), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1116), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1117), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n1118), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n1119), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n1120), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n1121), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n1122), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n1123), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n1124), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n1125), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n1126), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n1127), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n1128), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n1129), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n1130), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n1131), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n1132), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n1133), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n1134), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n1135), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n1136), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n1137), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n1138), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n1139), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n1140), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n1141), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n1142), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n1143), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n1144), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n1145), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n1146), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n1147), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n1148), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n1149), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n1150), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n1151), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n1152), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n1153), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n1154), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n1155), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n1156), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n1157), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n1158), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n1159), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n1160), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n1161), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n1162), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n1163), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n1164), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n1165), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n1166), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n1167), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n1168), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n1169), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n1170), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n1171), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n1172), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n1173), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n1174), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n1175), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n1176), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n1177), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n1178), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n1179), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n1180), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n1181), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n1182), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n1183), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n1184), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n1185), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n1186), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n1187), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n1188), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n1189), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n1190), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n1191), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n1192), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n1193), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n1194), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n1195), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n1196), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n1197), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n1198), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n1199), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n1200), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n1201), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n1202), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n1203), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n1204), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n1205), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n1206), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n1207), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n1208), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n1209), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n1210), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n1211), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n1212), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n1213), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n1214), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n1215), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n1216), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n1217), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n1218), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n1219), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n1220), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n1221), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n1222), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n1223), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n1224), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n1225), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n1226), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n1227), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n1228), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n1229), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n1230), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n1231), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n1232), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n1233), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n1234), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n1235), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n1236), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n1237), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n1238), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n1239), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n1240), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n1241), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n1242), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n1243), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n1244), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n1245), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n1246), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n1247), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n1248), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n1249), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n1250), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n1251), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n1252), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n1253), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n1254), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n1255), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n1256), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n1257), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n1258), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n1259), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n1260), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n1261), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n1262), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n1263), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n1264), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n1265), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n1266), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n1267), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n1268), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n1269), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n1270), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n1271), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n1272), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n1273), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n1274), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n1275), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n1276), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n1277), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n1278), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n1279), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n1280), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n1281), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n1282), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n1283), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n1284), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n1285), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n1286), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n1287), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n1288), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n1289), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n1290), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n1291), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n1292), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n1293), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n1294), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n1295), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n1296), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n1297), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n1298), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n1299), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n1300), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n1301), .CLK(clk), .Q(\mem<31><0> ) );
  DFFPOSX1 \mem_reg<32><7>  ( .D(n1302), .CLK(clk), .Q(\mem<32><7> ) );
  DFFPOSX1 \mem_reg<32><6>  ( .D(n1303), .CLK(clk), .Q(\mem<32><6> ) );
  DFFPOSX1 \mem_reg<32><5>  ( .D(n1304), .CLK(clk), .Q(\mem<32><5> ) );
  DFFPOSX1 \mem_reg<32><4>  ( .D(n1305), .CLK(clk), .Q(\mem<32><4> ) );
  DFFPOSX1 \mem_reg<32><3>  ( .D(n1306), .CLK(clk), .Q(\mem<32><3> ) );
  DFFPOSX1 \mem_reg<32><2>  ( .D(n1307), .CLK(clk), .Q(\mem<32><2> ) );
  DFFPOSX1 \mem_reg<32><1>  ( .D(n1308), .CLK(clk), .Q(\mem<32><1> ) );
  DFFPOSX1 \mem_reg<32><0>  ( .D(n1309), .CLK(clk), .Q(\mem<32><0> ) );
  AND2X2 U9 ( .A(n1477), .B(n1476), .Y(n1478) );
  AND2X2 U10 ( .A(n1472), .B(n1471), .Y(n1473) );
  AND2X2 U11 ( .A(n1466), .B(n1465), .Y(n1467) );
  AND2X2 U12 ( .A(n1461), .B(n1460), .Y(n1462) );
  AND2X2 U13 ( .A(n1455), .B(n1454), .Y(n1456) );
  AND2X2 U14 ( .A(n1450), .B(n1449), .Y(n1451) );
  AND2X2 U15 ( .A(n1444), .B(n1443), .Y(n1445) );
  AND2X2 U16 ( .A(n1439), .B(n1438), .Y(n1440) );
  AND2X2 U17 ( .A(n1433), .B(n1432), .Y(n1434) );
  AND2X2 U18 ( .A(n1428), .B(n1427), .Y(n1429) );
  AND2X2 U19 ( .A(n1422), .B(n1421), .Y(n1423) );
  AND2X2 U20 ( .A(n1417), .B(n1416), .Y(n1418) );
  AND2X2 U21 ( .A(n1411), .B(n1410), .Y(n1412) );
  AND2X2 U22 ( .A(n1406), .B(n1405), .Y(n1407) );
  AND2X2 U30 ( .A(n1326), .B(n1024), .Y(n1631) );
  AND2X2 U31 ( .A(n1325), .B(n1024), .Y(n1786) );
  AND2X2 U32 ( .A(n1326), .B(\addr_1c<0> ), .Y(n1651) );
  AND2X2 U33 ( .A(n1325), .B(\addr_1c<0> ), .Y(n1806) );
  AND2X2 U34 ( .A(n1320), .B(n1319), .Y(n1321) );
  AND2X2 U45 ( .A(n1313), .B(n1312), .Y(n1314) );
  NOR3X1 U94 ( .A(n1044), .B(rd), .C(n963), .Y(wr0) );
  NOR3X1 U95 ( .A(n1045), .B(wr), .C(n963), .Y(rd0) );
  OAI21X1 U96 ( .A(n1011), .B(n1036), .C(n1836), .Y(n1309) );
  NAND2X1 U97 ( .A(\mem<32><0> ), .B(n1011), .Y(n1836) );
  OAI21X1 U98 ( .A(n1011), .B(n1037), .C(n1835), .Y(n1308) );
  NAND2X1 U99 ( .A(\mem<32><1> ), .B(n1011), .Y(n1835) );
  OAI21X1 U100 ( .A(n1011), .B(n1038), .C(n1834), .Y(n1307) );
  NAND2X1 U101 ( .A(\mem<32><2> ), .B(n1011), .Y(n1834) );
  OAI21X1 U102 ( .A(n1011), .B(n1039), .C(n1833), .Y(n1306) );
  NAND2X1 U103 ( .A(\mem<32><3> ), .B(n1011), .Y(n1833) );
  OAI21X1 U104 ( .A(n1011), .B(n1040), .C(n1832), .Y(n1305) );
  NAND2X1 U105 ( .A(\mem<32><4> ), .B(n1011), .Y(n1832) );
  OAI21X1 U106 ( .A(n1011), .B(n1041), .C(n1831), .Y(n1304) );
  NAND2X1 U107 ( .A(\mem<32><5> ), .B(n1011), .Y(n1831) );
  OAI21X1 U108 ( .A(n1011), .B(n1042), .C(n1830), .Y(n1303) );
  NAND2X1 U109 ( .A(\mem<32><6> ), .B(n1011), .Y(n1830) );
  OAI21X1 U110 ( .A(n1011), .B(n1043), .C(n1829), .Y(n1302) );
  NAND2X1 U111 ( .A(\mem<32><7> ), .B(n1011), .Y(n1829) );
  NAND3X1 U112 ( .A(n1828), .B(n1827), .C(n964), .Y(n1837) );
  OAI21X1 U113 ( .A(n6), .B(n1028), .C(n1826), .Y(n1301) );
  NAND2X1 U114 ( .A(\mem<31><0> ), .B(n6), .Y(n1826) );
  OAI21X1 U115 ( .A(n6), .B(n1029), .C(n1825), .Y(n1300) );
  NAND2X1 U116 ( .A(\mem<31><1> ), .B(n6), .Y(n1825) );
  OAI21X1 U117 ( .A(n6), .B(n1030), .C(n1824), .Y(n1299) );
  NAND2X1 U118 ( .A(\mem<31><2> ), .B(n6), .Y(n1824) );
  OAI21X1 U119 ( .A(n6), .B(n1031), .C(n1823), .Y(n1298) );
  NAND2X1 U120 ( .A(\mem<31><3> ), .B(n6), .Y(n1823) );
  OAI21X1 U121 ( .A(n6), .B(n1032), .C(n1822), .Y(n1297) );
  NAND2X1 U122 ( .A(\mem<31><4> ), .B(n6), .Y(n1822) );
  OAI21X1 U123 ( .A(n6), .B(n1033), .C(n1821), .Y(n1296) );
  NAND2X1 U124 ( .A(\mem<31><5> ), .B(n6), .Y(n1821) );
  OAI21X1 U125 ( .A(n6), .B(n1034), .C(n1820), .Y(n1295) );
  NAND2X1 U126 ( .A(\mem<31><6> ), .B(n6), .Y(n1820) );
  OAI21X1 U127 ( .A(n6), .B(n1035), .C(n1819), .Y(n1294) );
  NAND2X1 U128 ( .A(\mem<31><7> ), .B(n6), .Y(n1819) );
  OAI21X1 U130 ( .A(n1036), .B(n1010), .C(n1815), .Y(n1293) );
  NAND2X1 U131 ( .A(\mem<30><0> ), .B(n1010), .Y(n1815) );
  OAI21X1 U132 ( .A(n1037), .B(n1009), .C(n1814), .Y(n1292) );
  NAND2X1 U133 ( .A(\mem<30><1> ), .B(n1010), .Y(n1814) );
  OAI21X1 U134 ( .A(n1038), .B(n1009), .C(n1813), .Y(n1291) );
  NAND2X1 U135 ( .A(\mem<30><2> ), .B(n1010), .Y(n1813) );
  OAI21X1 U136 ( .A(n1039), .B(n1009), .C(n1812), .Y(n1290) );
  NAND2X1 U137 ( .A(\mem<30><3> ), .B(n1010), .Y(n1812) );
  OAI21X1 U138 ( .A(n1040), .B(n1009), .C(n1811), .Y(n1289) );
  NAND2X1 U139 ( .A(\mem<30><4> ), .B(n1010), .Y(n1811) );
  OAI21X1 U140 ( .A(n1041), .B(n1009), .C(n1810), .Y(n1288) );
  NAND2X1 U141 ( .A(\mem<30><5> ), .B(n1010), .Y(n1810) );
  OAI21X1 U142 ( .A(n1042), .B(n1009), .C(n1809), .Y(n1287) );
  NAND2X1 U143 ( .A(\mem<30><6> ), .B(n1010), .Y(n1809) );
  OAI21X1 U144 ( .A(n1043), .B(n1009), .C(n1808), .Y(n1286) );
  NAND2X1 U145 ( .A(\mem<30><7> ), .B(n1010), .Y(n1808) );
  NAND3X1 U146 ( .A(n1807), .B(n1828), .C(n1806), .Y(n1816) );
  OAI21X1 U147 ( .A(n1028), .B(n1008), .C(n1804), .Y(n1285) );
  NAND2X1 U148 ( .A(\mem<29><0> ), .B(n1008), .Y(n1804) );
  OAI21X1 U149 ( .A(n1029), .B(n1008), .C(n1803), .Y(n1284) );
  NAND2X1 U150 ( .A(\mem<29><1> ), .B(n1008), .Y(n1803) );
  OAI21X1 U151 ( .A(n1030), .B(n1008), .C(n1802), .Y(n1283) );
  NAND2X1 U152 ( .A(\mem<29><2> ), .B(n1008), .Y(n1802) );
  OAI21X1 U153 ( .A(n1031), .B(n1008), .C(n1801), .Y(n1282) );
  NAND2X1 U154 ( .A(\mem<29><3> ), .B(n1008), .Y(n1801) );
  OAI21X1 U155 ( .A(n1032), .B(n1008), .C(n1800), .Y(n1281) );
  NAND2X1 U156 ( .A(\mem<29><4> ), .B(n1008), .Y(n1800) );
  OAI21X1 U157 ( .A(n1033), .B(n1008), .C(n1799), .Y(n1280) );
  NAND2X1 U158 ( .A(\mem<29><5> ), .B(n1008), .Y(n1799) );
  OAI21X1 U159 ( .A(n1034), .B(n1008), .C(n1798), .Y(n1279) );
  NAND2X1 U160 ( .A(\mem<29><6> ), .B(n1008), .Y(n1798) );
  OAI21X1 U161 ( .A(n1035), .B(n1008), .C(n1797), .Y(n1278) );
  NAND2X1 U162 ( .A(\mem<29><7> ), .B(n1008), .Y(n1797) );
  NAND3X1 U163 ( .A(n973), .B(n1828), .C(n1796), .Y(n1805) );
  OAI21X1 U164 ( .A(n1036), .B(n1007), .C(n1794), .Y(n1277) );
  NAND2X1 U165 ( .A(\mem<28><0> ), .B(n1007), .Y(n1794) );
  OAI21X1 U166 ( .A(n1037), .B(n1006), .C(n1793), .Y(n1276) );
  NAND2X1 U167 ( .A(\mem<28><1> ), .B(n1007), .Y(n1793) );
  OAI21X1 U168 ( .A(n1038), .B(n1006), .C(n1792), .Y(n1275) );
  NAND2X1 U169 ( .A(\mem<28><2> ), .B(n1007), .Y(n1792) );
  OAI21X1 U170 ( .A(n1039), .B(n1006), .C(n1791), .Y(n1274) );
  NAND2X1 U171 ( .A(\mem<28><3> ), .B(n1007), .Y(n1791) );
  OAI21X1 U172 ( .A(n1040), .B(n1006), .C(n1790), .Y(n1273) );
  NAND2X1 U173 ( .A(\mem<28><4> ), .B(n1007), .Y(n1790) );
  OAI21X1 U174 ( .A(n1041), .B(n1006), .C(n1789), .Y(n1272) );
  NAND2X1 U175 ( .A(\mem<28><5> ), .B(n1007), .Y(n1789) );
  OAI21X1 U176 ( .A(n1042), .B(n1006), .C(n1788), .Y(n1271) );
  NAND2X1 U177 ( .A(\mem<28><6> ), .B(n1007), .Y(n1788) );
  OAI21X1 U178 ( .A(n1043), .B(n1006), .C(n1787), .Y(n1270) );
  NAND2X1 U179 ( .A(\mem<28><7> ), .B(n1007), .Y(n1787) );
  NAND3X1 U180 ( .A(n1807), .B(n1828), .C(n1786), .Y(n1795) );
  OAI21X1 U181 ( .A(n1028), .B(n1005), .C(n1784), .Y(n1269) );
  NAND2X1 U182 ( .A(\mem<27><0> ), .B(n1005), .Y(n1784) );
  OAI21X1 U183 ( .A(n1029), .B(n1005), .C(n1783), .Y(n1268) );
  NAND2X1 U184 ( .A(\mem<27><1> ), .B(n1005), .Y(n1783) );
  OAI21X1 U185 ( .A(n1030), .B(n1005), .C(n1782), .Y(n1267) );
  NAND2X1 U186 ( .A(\mem<27><2> ), .B(n1005), .Y(n1782) );
  OAI21X1 U187 ( .A(n1031), .B(n1005), .C(n1781), .Y(n1266) );
  NAND2X1 U188 ( .A(\mem<27><3> ), .B(n1005), .Y(n1781) );
  OAI21X1 U189 ( .A(n1032), .B(n1005), .C(n1780), .Y(n1265) );
  NAND2X1 U190 ( .A(\mem<27><4> ), .B(n1005), .Y(n1780) );
  OAI21X1 U191 ( .A(n1033), .B(n1005), .C(n1779), .Y(n1264) );
  NAND2X1 U192 ( .A(\mem<27><5> ), .B(n1005), .Y(n1779) );
  OAI21X1 U193 ( .A(n1034), .B(n1005), .C(n1778), .Y(n1263) );
  NAND2X1 U194 ( .A(\mem<27><6> ), .B(n1005), .Y(n1778) );
  OAI21X1 U195 ( .A(n1035), .B(n1005), .C(n1777), .Y(n1262) );
  NAND2X1 U196 ( .A(\mem<27><7> ), .B(n1005), .Y(n1777) );
  NAND3X1 U197 ( .A(n973), .B(n1828), .C(n1776), .Y(n1785) );
  OAI21X1 U198 ( .A(n1036), .B(n1004), .C(n1774), .Y(n1261) );
  NAND2X1 U199 ( .A(\mem<26><0> ), .B(n1004), .Y(n1774) );
  OAI21X1 U200 ( .A(n1037), .B(n1003), .C(n1773), .Y(n1260) );
  NAND2X1 U201 ( .A(\mem<26><1> ), .B(n1004), .Y(n1773) );
  OAI21X1 U202 ( .A(n1038), .B(n1003), .C(n1772), .Y(n1259) );
  NAND2X1 U203 ( .A(\mem<26><2> ), .B(n1004), .Y(n1772) );
  OAI21X1 U204 ( .A(n1039), .B(n1003), .C(n1771), .Y(n1258) );
  NAND2X1 U205 ( .A(\mem<26><3> ), .B(n1004), .Y(n1771) );
  OAI21X1 U206 ( .A(n1040), .B(n1003), .C(n1770), .Y(n1257) );
  NAND2X1 U207 ( .A(\mem<26><4> ), .B(n1004), .Y(n1770) );
  OAI21X1 U208 ( .A(n1041), .B(n1003), .C(n1769), .Y(n1256) );
  NAND2X1 U209 ( .A(\mem<26><5> ), .B(n1004), .Y(n1769) );
  OAI21X1 U210 ( .A(n1042), .B(n1003), .C(n1768), .Y(n1255) );
  NAND2X1 U211 ( .A(\mem<26><6> ), .B(n1004), .Y(n1768) );
  OAI21X1 U212 ( .A(n1043), .B(n1003), .C(n1767), .Y(n1254) );
  NAND2X1 U213 ( .A(\mem<26><7> ), .B(n1004), .Y(n1767) );
  NAND3X1 U214 ( .A(n1806), .B(n1828), .C(n1766), .Y(n1775) );
  OAI21X1 U215 ( .A(n1028), .B(n1002), .C(n1764), .Y(n1253) );
  NAND2X1 U216 ( .A(\mem<25><0> ), .B(n1002), .Y(n1764) );
  OAI21X1 U217 ( .A(n1029), .B(n1002), .C(n1763), .Y(n1252) );
  NAND2X1 U218 ( .A(\mem<25><1> ), .B(n1002), .Y(n1763) );
  OAI21X1 U219 ( .A(n1030), .B(n1002), .C(n1762), .Y(n1251) );
  NAND2X1 U220 ( .A(\mem<25><2> ), .B(n1002), .Y(n1762) );
  OAI21X1 U221 ( .A(n1031), .B(n1002), .C(n1761), .Y(n1250) );
  NAND2X1 U222 ( .A(\mem<25><3> ), .B(n1002), .Y(n1761) );
  OAI21X1 U223 ( .A(n1032), .B(n1002), .C(n1760), .Y(n1249) );
  NAND2X1 U224 ( .A(\mem<25><4> ), .B(n1002), .Y(n1760) );
  OAI21X1 U225 ( .A(n1033), .B(n1002), .C(n1759), .Y(n1248) );
  NAND2X1 U226 ( .A(\mem<25><5> ), .B(n1002), .Y(n1759) );
  OAI21X1 U227 ( .A(n1034), .B(n1002), .C(n1758), .Y(n1247) );
  NAND2X1 U228 ( .A(\mem<25><6> ), .B(n1002), .Y(n1758) );
  OAI21X1 U229 ( .A(n1035), .B(n1002), .C(n1757), .Y(n1246) );
  NAND2X1 U230 ( .A(\mem<25><7> ), .B(n1002), .Y(n1757) );
  NAND3X1 U231 ( .A(n973), .B(n1828), .C(n1756), .Y(n1765) );
  OAI21X1 U232 ( .A(n1036), .B(n1001), .C(n1754), .Y(n1245) );
  NAND2X1 U233 ( .A(\mem<24><0> ), .B(n1001), .Y(n1754) );
  OAI21X1 U234 ( .A(n1037), .B(n1000), .C(n1753), .Y(n1244) );
  NAND2X1 U235 ( .A(\mem<24><1> ), .B(n1001), .Y(n1753) );
  OAI21X1 U236 ( .A(n1038), .B(n1000), .C(n1752), .Y(n1243) );
  NAND2X1 U237 ( .A(\mem<24><2> ), .B(n1001), .Y(n1752) );
  OAI21X1 U238 ( .A(n1039), .B(n1000), .C(n1751), .Y(n1242) );
  NAND2X1 U239 ( .A(\mem<24><3> ), .B(n1001), .Y(n1751) );
  OAI21X1 U240 ( .A(n1040), .B(n1000), .C(n1750), .Y(n1241) );
  NAND2X1 U241 ( .A(\mem<24><4> ), .B(n1001), .Y(n1750) );
  OAI21X1 U242 ( .A(n1041), .B(n1000), .C(n1749), .Y(n1240) );
  NAND2X1 U243 ( .A(\mem<24><5> ), .B(n1001), .Y(n1749) );
  OAI21X1 U244 ( .A(n1042), .B(n1000), .C(n1748), .Y(n1239) );
  NAND2X1 U245 ( .A(\mem<24><6> ), .B(n1001), .Y(n1748) );
  OAI21X1 U246 ( .A(n1043), .B(n1000), .C(n1747), .Y(n1238) );
  NAND2X1 U247 ( .A(\mem<24><7> ), .B(n1001), .Y(n1747) );
  NAND3X1 U248 ( .A(n1786), .B(n1828), .C(n1766), .Y(n1755) );
  OAI21X1 U249 ( .A(n1028), .B(n999), .C(n1745), .Y(n1237) );
  NAND2X1 U250 ( .A(\mem<23><0> ), .B(n999), .Y(n1745) );
  OAI21X1 U251 ( .A(n1029), .B(n999), .C(n1744), .Y(n1236) );
  NAND2X1 U252 ( .A(\mem<23><1> ), .B(n999), .Y(n1744) );
  OAI21X1 U253 ( .A(n1030), .B(n999), .C(n1743), .Y(n1235) );
  NAND2X1 U254 ( .A(\mem<23><2> ), .B(n999), .Y(n1743) );
  OAI21X1 U255 ( .A(n1031), .B(n999), .C(n1742), .Y(n1234) );
  NAND2X1 U256 ( .A(\mem<23><3> ), .B(n999), .Y(n1742) );
  OAI21X1 U257 ( .A(n1032), .B(n999), .C(n1741), .Y(n1233) );
  NAND2X1 U258 ( .A(\mem<23><4> ), .B(n999), .Y(n1741) );
  OAI21X1 U259 ( .A(n1033), .B(n999), .C(n1740), .Y(n1232) );
  NAND2X1 U260 ( .A(\mem<23><5> ), .B(n999), .Y(n1740) );
  OAI21X1 U261 ( .A(n1034), .B(n999), .C(n1739), .Y(n1231) );
  NAND2X1 U262 ( .A(\mem<23><6> ), .B(n999), .Y(n1739) );
  OAI21X1 U263 ( .A(n1035), .B(n999), .C(n1738), .Y(n1230) );
  NAND2X1 U264 ( .A(\mem<23><7> ), .B(n999), .Y(n1738) );
  NAND3X1 U265 ( .A(n973), .B(n1828), .C(n1737), .Y(n1746) );
  OAI21X1 U266 ( .A(n1036), .B(n998), .C(n1735), .Y(n1229) );
  NAND2X1 U267 ( .A(\mem<22><0> ), .B(n998), .Y(n1735) );
  OAI21X1 U268 ( .A(n1037), .B(n998), .C(n1734), .Y(n1228) );
  NAND2X1 U269 ( .A(\mem<22><1> ), .B(n998), .Y(n1734) );
  OAI21X1 U270 ( .A(n1038), .B(n998), .C(n1733), .Y(n1227) );
  NAND2X1 U271 ( .A(\mem<22><2> ), .B(n998), .Y(n1733) );
  OAI21X1 U272 ( .A(n1039), .B(n998), .C(n1732), .Y(n1226) );
  NAND2X1 U273 ( .A(\mem<22><3> ), .B(n998), .Y(n1732) );
  OAI21X1 U274 ( .A(n1040), .B(n998), .C(n1731), .Y(n1225) );
  NAND2X1 U275 ( .A(\mem<22><4> ), .B(n998), .Y(n1731) );
  OAI21X1 U276 ( .A(n1041), .B(n998), .C(n1730), .Y(n1224) );
  NAND2X1 U277 ( .A(\mem<22><5> ), .B(n998), .Y(n1730) );
  OAI21X1 U278 ( .A(n1042), .B(n998), .C(n1729), .Y(n1223) );
  NAND2X1 U279 ( .A(\mem<22><6> ), .B(n998), .Y(n1729) );
  OAI21X1 U280 ( .A(n1043), .B(n998), .C(n1728), .Y(n1222) );
  NAND2X1 U281 ( .A(\mem<22><7> ), .B(n998), .Y(n1728) );
  NAND3X1 U282 ( .A(n1806), .B(n1828), .C(n969), .Y(n1736) );
  OAI21X1 U283 ( .A(n1028), .B(n997), .C(n1726), .Y(n1221) );
  NAND2X1 U284 ( .A(\mem<21><0> ), .B(n997), .Y(n1726) );
  OAI21X1 U285 ( .A(n1029), .B(n997), .C(n1725), .Y(n1220) );
  NAND2X1 U286 ( .A(\mem<21><1> ), .B(n997), .Y(n1725) );
  OAI21X1 U287 ( .A(n1030), .B(n997), .C(n1724), .Y(n1219) );
  NAND2X1 U288 ( .A(\mem<21><2> ), .B(n997), .Y(n1724) );
  OAI21X1 U289 ( .A(n1031), .B(n997), .C(n1723), .Y(n1218) );
  NAND2X1 U290 ( .A(\mem<21><3> ), .B(n997), .Y(n1723) );
  OAI21X1 U291 ( .A(n1032), .B(n997), .C(n1722), .Y(n1217) );
  NAND2X1 U292 ( .A(\mem<21><4> ), .B(n997), .Y(n1722) );
  OAI21X1 U293 ( .A(n1033), .B(n997), .C(n1721), .Y(n1216) );
  NAND2X1 U294 ( .A(\mem<21><5> ), .B(n997), .Y(n1721) );
  OAI21X1 U295 ( .A(n1034), .B(n997), .C(n1720), .Y(n1215) );
  NAND2X1 U296 ( .A(\mem<21><6> ), .B(n997), .Y(n1720) );
  OAI21X1 U297 ( .A(n1035), .B(n997), .C(n1719), .Y(n1214) );
  NAND2X1 U298 ( .A(\mem<21><7> ), .B(n997), .Y(n1719) );
  NAND3X1 U299 ( .A(n973), .B(n1828), .C(n1718), .Y(n1727) );
  OAI21X1 U300 ( .A(n1036), .B(n996), .C(n1716), .Y(n1213) );
  NAND2X1 U301 ( .A(\mem<20><0> ), .B(n996), .Y(n1716) );
  OAI21X1 U302 ( .A(n1037), .B(n996), .C(n1715), .Y(n1212) );
  NAND2X1 U303 ( .A(\mem<20><1> ), .B(n996), .Y(n1715) );
  OAI21X1 U304 ( .A(n1038), .B(n996), .C(n1714), .Y(n1211) );
  NAND2X1 U305 ( .A(\mem<20><2> ), .B(n996), .Y(n1714) );
  OAI21X1 U306 ( .A(n1039), .B(n996), .C(n1713), .Y(n1210) );
  NAND2X1 U307 ( .A(\mem<20><3> ), .B(n996), .Y(n1713) );
  OAI21X1 U308 ( .A(n1040), .B(n996), .C(n1712), .Y(n1209) );
  NAND2X1 U309 ( .A(\mem<20><4> ), .B(n996), .Y(n1712) );
  OAI21X1 U310 ( .A(n1041), .B(n996), .C(n1711), .Y(n1208) );
  NAND2X1 U311 ( .A(\mem<20><5> ), .B(n996), .Y(n1711) );
  OAI21X1 U312 ( .A(n1042), .B(n996), .C(n1710), .Y(n1207) );
  NAND2X1 U313 ( .A(\mem<20><6> ), .B(n996), .Y(n1710) );
  OAI21X1 U314 ( .A(n1043), .B(n996), .C(n1709), .Y(n1206) );
  NAND2X1 U315 ( .A(\mem<20><7> ), .B(n996), .Y(n1709) );
  NAND3X1 U316 ( .A(n1786), .B(n1828), .C(n969), .Y(n1717) );
  OAI21X1 U317 ( .A(n1028), .B(n995), .C(n1707), .Y(n1205) );
  NAND2X1 U318 ( .A(\mem<19><0> ), .B(n995), .Y(n1707) );
  OAI21X1 U319 ( .A(n1029), .B(n995), .C(n1706), .Y(n1204) );
  NAND2X1 U320 ( .A(\mem<19><1> ), .B(n995), .Y(n1706) );
  OAI21X1 U321 ( .A(n1030), .B(n995), .C(n1705), .Y(n1203) );
  NAND2X1 U322 ( .A(\mem<19><2> ), .B(n995), .Y(n1705) );
  OAI21X1 U323 ( .A(n1031), .B(n995), .C(n1704), .Y(n1202) );
  NAND2X1 U324 ( .A(\mem<19><3> ), .B(n995), .Y(n1704) );
  OAI21X1 U325 ( .A(n1032), .B(n995), .C(n1703), .Y(n1201) );
  NAND2X1 U326 ( .A(\mem<19><4> ), .B(n995), .Y(n1703) );
  OAI21X1 U327 ( .A(n1033), .B(n995), .C(n1702), .Y(n1200) );
  NAND2X1 U328 ( .A(\mem<19><5> ), .B(n995), .Y(n1702) );
  OAI21X1 U329 ( .A(n1034), .B(n995), .C(n1701), .Y(n1199) );
  NAND2X1 U330 ( .A(\mem<19><6> ), .B(n995), .Y(n1701) );
  OAI21X1 U331 ( .A(n1035), .B(n995), .C(n1700), .Y(n1198) );
  NAND2X1 U332 ( .A(\mem<19><7> ), .B(n995), .Y(n1700) );
  NAND3X1 U333 ( .A(n973), .B(n1828), .C(n1699), .Y(n1708) );
  OAI21X1 U334 ( .A(n1036), .B(n994), .C(n1697), .Y(n1197) );
  NAND2X1 U335 ( .A(\mem<18><0> ), .B(n994), .Y(n1697) );
  OAI21X1 U336 ( .A(n1037), .B(n994), .C(n1696), .Y(n1196) );
  NAND2X1 U337 ( .A(\mem<18><1> ), .B(n994), .Y(n1696) );
  OAI21X1 U338 ( .A(n1038), .B(n994), .C(n1695), .Y(n1195) );
  NAND2X1 U339 ( .A(\mem<18><2> ), .B(n994), .Y(n1695) );
  OAI21X1 U340 ( .A(n1039), .B(n994), .C(n1694), .Y(n1194) );
  NAND2X1 U341 ( .A(\mem<18><3> ), .B(n994), .Y(n1694) );
  OAI21X1 U342 ( .A(n1040), .B(n994), .C(n1693), .Y(n1193) );
  NAND2X1 U343 ( .A(\mem<18><4> ), .B(n994), .Y(n1693) );
  OAI21X1 U344 ( .A(n1041), .B(n994), .C(n1692), .Y(n1192) );
  NAND2X1 U345 ( .A(\mem<18><5> ), .B(n994), .Y(n1692) );
  OAI21X1 U346 ( .A(n1042), .B(n994), .C(n1691), .Y(n1191) );
  NAND2X1 U347 ( .A(\mem<18><6> ), .B(n994), .Y(n1691) );
  OAI21X1 U348 ( .A(n1043), .B(n994), .C(n1690), .Y(n1190) );
  NAND2X1 U349 ( .A(\mem<18><7> ), .B(n994), .Y(n1690) );
  NAND3X1 U350 ( .A(n1806), .B(n1828), .C(n967), .Y(n1698) );
  OAI21X1 U351 ( .A(n1028), .B(n993), .C(n1688), .Y(n1189) );
  NAND2X1 U352 ( .A(\mem<17><0> ), .B(n993), .Y(n1688) );
  OAI21X1 U353 ( .A(n1029), .B(n993), .C(n1687), .Y(n1188) );
  NAND2X1 U354 ( .A(\mem<17><1> ), .B(n993), .Y(n1687) );
  OAI21X1 U355 ( .A(n1030), .B(n993), .C(n1686), .Y(n1187) );
  NAND2X1 U356 ( .A(\mem<17><2> ), .B(n993), .Y(n1686) );
  OAI21X1 U357 ( .A(n1031), .B(n993), .C(n1685), .Y(n1186) );
  NAND2X1 U358 ( .A(\mem<17><3> ), .B(n993), .Y(n1685) );
  OAI21X1 U359 ( .A(n1032), .B(n993), .C(n1684), .Y(n1185) );
  NAND2X1 U360 ( .A(\mem<17><4> ), .B(n993), .Y(n1684) );
  OAI21X1 U361 ( .A(n1033), .B(n993), .C(n1683), .Y(n1184) );
  NAND2X1 U362 ( .A(\mem<17><5> ), .B(n993), .Y(n1683) );
  OAI21X1 U363 ( .A(n1034), .B(n993), .C(n1682), .Y(n1183) );
  NAND2X1 U364 ( .A(\mem<17><6> ), .B(n993), .Y(n1682) );
  OAI21X1 U365 ( .A(n1035), .B(n993), .C(n1681), .Y(n1182) );
  NAND2X1 U366 ( .A(\mem<17><7> ), .B(n993), .Y(n1681) );
  NAND3X1 U367 ( .A(n973), .B(n1828), .C(n1680), .Y(n1689) );
  OAI21X1 U368 ( .A(n1036), .B(n992), .C(n1678), .Y(n1181) );
  NAND2X1 U369 ( .A(\mem<16><0> ), .B(n992), .Y(n1678) );
  OAI21X1 U370 ( .A(n1037), .B(n992), .C(n1677), .Y(n1180) );
  NAND2X1 U371 ( .A(\mem<16><1> ), .B(n992), .Y(n1677) );
  OAI21X1 U372 ( .A(n1038), .B(n992), .C(n1676), .Y(n1179) );
  NAND2X1 U373 ( .A(\mem<16><2> ), .B(n992), .Y(n1676) );
  OAI21X1 U374 ( .A(n1039), .B(n992), .C(n1675), .Y(n1178) );
  NAND2X1 U375 ( .A(\mem<16><3> ), .B(n992), .Y(n1675) );
  OAI21X1 U376 ( .A(n1040), .B(n992), .C(n1674), .Y(n1177) );
  NAND2X1 U377 ( .A(\mem<16><4> ), .B(n992), .Y(n1674) );
  OAI21X1 U378 ( .A(n1041), .B(n992), .C(n1673), .Y(n1176) );
  NAND2X1 U379 ( .A(\mem<16><5> ), .B(n992), .Y(n1673) );
  OAI21X1 U380 ( .A(n1042), .B(n992), .C(n1672), .Y(n1175) );
  NAND2X1 U381 ( .A(\mem<16><6> ), .B(n992), .Y(n1672) );
  OAI21X1 U382 ( .A(n1043), .B(n992), .C(n1671), .Y(n1174) );
  NAND2X1 U383 ( .A(\mem<16><7> ), .B(n992), .Y(n1671) );
  NAND3X1 U384 ( .A(n1786), .B(n1828), .C(n967), .Y(n1679) );
  OAI21X1 U385 ( .A(n1028), .B(n991), .C(n1669), .Y(n1173) );
  NAND2X1 U386 ( .A(\mem<15><0> ), .B(n991), .Y(n1669) );
  OAI21X1 U387 ( .A(n1029), .B(n991), .C(n1668), .Y(n1172) );
  NAND2X1 U388 ( .A(\mem<15><1> ), .B(n991), .Y(n1668) );
  OAI21X1 U389 ( .A(n1030), .B(n991), .C(n1667), .Y(n1171) );
  NAND2X1 U390 ( .A(\mem<15><2> ), .B(n991), .Y(n1667) );
  OAI21X1 U391 ( .A(n1031), .B(n991), .C(n1666), .Y(n1170) );
  NAND2X1 U392 ( .A(\mem<15><3> ), .B(n991), .Y(n1666) );
  OAI21X1 U393 ( .A(n1032), .B(n991), .C(n1665), .Y(n1169) );
  NAND2X1 U394 ( .A(\mem<15><4> ), .B(n991), .Y(n1665) );
  OAI21X1 U395 ( .A(n1033), .B(n991), .C(n1664), .Y(n1168) );
  NAND2X1 U396 ( .A(\mem<15><5> ), .B(n991), .Y(n1664) );
  OAI21X1 U397 ( .A(n1034), .B(n991), .C(n1663), .Y(n1167) );
  NAND2X1 U398 ( .A(\mem<15><6> ), .B(n991), .Y(n1663) );
  OAI21X1 U399 ( .A(n1035), .B(n991), .C(n1662), .Y(n1166) );
  NAND2X1 U400 ( .A(\mem<15><7> ), .B(n991), .Y(n1662) );
  NAND3X1 U401 ( .A(n973), .B(n1828), .C(n1661), .Y(n1670) );
  OAI21X1 U402 ( .A(n1036), .B(n990), .C(n1659), .Y(n1165) );
  NAND2X1 U403 ( .A(\mem<14><0> ), .B(n990), .Y(n1659) );
  OAI21X1 U404 ( .A(n1037), .B(n989), .C(n1658), .Y(n1164) );
  NAND2X1 U405 ( .A(\mem<14><1> ), .B(n990), .Y(n1658) );
  OAI21X1 U406 ( .A(n1038), .B(n989), .C(n1657), .Y(n1163) );
  NAND2X1 U407 ( .A(\mem<14><2> ), .B(n990), .Y(n1657) );
  OAI21X1 U408 ( .A(n1039), .B(n989), .C(n1656), .Y(n1162) );
  NAND2X1 U409 ( .A(\mem<14><3> ), .B(n990), .Y(n1656) );
  OAI21X1 U410 ( .A(n1040), .B(n989), .C(n1655), .Y(n1161) );
  NAND2X1 U411 ( .A(\mem<14><4> ), .B(n990), .Y(n1655) );
  OAI21X1 U412 ( .A(n1041), .B(n989), .C(n1654), .Y(n1160) );
  NAND2X1 U413 ( .A(\mem<14><5> ), .B(n990), .Y(n1654) );
  OAI21X1 U414 ( .A(n1042), .B(n989), .C(n1653), .Y(n1159) );
  NAND2X1 U415 ( .A(\mem<14><6> ), .B(n990), .Y(n1653) );
  OAI21X1 U416 ( .A(n1043), .B(n989), .C(n1652), .Y(n1158) );
  NAND2X1 U417 ( .A(\mem<14><7> ), .B(n990), .Y(n1652) );
  NAND3X1 U418 ( .A(n1807), .B(n1828), .C(n1651), .Y(n1660) );
  OAI21X1 U419 ( .A(n1028), .B(n988), .C(n1649), .Y(n1157) );
  NAND2X1 U420 ( .A(\mem<13><0> ), .B(n988), .Y(n1649) );
  OAI21X1 U421 ( .A(n1029), .B(n988), .C(n1648), .Y(n1156) );
  NAND2X1 U422 ( .A(\mem<13><1> ), .B(n988), .Y(n1648) );
  OAI21X1 U423 ( .A(n1030), .B(n988), .C(n1647), .Y(n1155) );
  NAND2X1 U424 ( .A(\mem<13><2> ), .B(n988), .Y(n1647) );
  OAI21X1 U425 ( .A(n1031), .B(n988), .C(n1646), .Y(n1154) );
  NAND2X1 U426 ( .A(\mem<13><3> ), .B(n988), .Y(n1646) );
  OAI21X1 U427 ( .A(n1032), .B(n988), .C(n1645), .Y(n1153) );
  NAND2X1 U428 ( .A(\mem<13><4> ), .B(n988), .Y(n1645) );
  OAI21X1 U429 ( .A(n1033), .B(n988), .C(n1644), .Y(n1152) );
  NAND2X1 U430 ( .A(\mem<13><5> ), .B(n988), .Y(n1644) );
  OAI21X1 U431 ( .A(n1034), .B(n988), .C(n1643), .Y(n1151) );
  NAND2X1 U432 ( .A(\mem<13><6> ), .B(n988), .Y(n1643) );
  OAI21X1 U433 ( .A(n1035), .B(n988), .C(n1642), .Y(n1150) );
  NAND2X1 U434 ( .A(\mem<13><7> ), .B(n988), .Y(n1642) );
  NAND3X1 U435 ( .A(n973), .B(n1828), .C(n1641), .Y(n1650) );
  OAI21X1 U436 ( .A(n1036), .B(n987), .C(n1639), .Y(n1149) );
  NAND2X1 U437 ( .A(\mem<12><0> ), .B(n987), .Y(n1639) );
  OAI21X1 U438 ( .A(n1037), .B(n986), .C(n1638), .Y(n1148) );
  NAND2X1 U439 ( .A(\mem<12><1> ), .B(n987), .Y(n1638) );
  OAI21X1 U440 ( .A(n1038), .B(n986), .C(n1637), .Y(n1147) );
  NAND2X1 U441 ( .A(\mem<12><2> ), .B(n987), .Y(n1637) );
  OAI21X1 U442 ( .A(n1039), .B(n986), .C(n1636), .Y(n1146) );
  NAND2X1 U443 ( .A(\mem<12><3> ), .B(n987), .Y(n1636) );
  OAI21X1 U444 ( .A(n1040), .B(n986), .C(n1635), .Y(n1145) );
  NAND2X1 U445 ( .A(\mem<12><4> ), .B(n987), .Y(n1635) );
  OAI21X1 U446 ( .A(n1041), .B(n986), .C(n1634), .Y(n1144) );
  NAND2X1 U447 ( .A(\mem<12><5> ), .B(n987), .Y(n1634) );
  OAI21X1 U448 ( .A(n1042), .B(n986), .C(n1633), .Y(n1143) );
  NAND2X1 U449 ( .A(\mem<12><6> ), .B(n987), .Y(n1633) );
  OAI21X1 U450 ( .A(n1043), .B(n986), .C(n1632), .Y(n1142) );
  NAND2X1 U451 ( .A(\mem<12><7> ), .B(n987), .Y(n1632) );
  NAND3X1 U452 ( .A(n1807), .B(n1828), .C(n1631), .Y(n1640) );
  OAI21X1 U453 ( .A(n1028), .B(n985), .C(n1628), .Y(n1141) );
  NAND2X1 U454 ( .A(\mem<11><0> ), .B(n985), .Y(n1628) );
  OAI21X1 U455 ( .A(n1029), .B(n985), .C(n1627), .Y(n1140) );
  NAND2X1 U456 ( .A(\mem<11><1> ), .B(n985), .Y(n1627) );
  OAI21X1 U457 ( .A(n1030), .B(n985), .C(n1626), .Y(n1139) );
  NAND2X1 U458 ( .A(\mem<11><2> ), .B(n985), .Y(n1626) );
  OAI21X1 U459 ( .A(n1031), .B(n985), .C(n1625), .Y(n1138) );
  NAND2X1 U460 ( .A(\mem<11><3> ), .B(n985), .Y(n1625) );
  OAI21X1 U461 ( .A(n1032), .B(n985), .C(n1624), .Y(n1137) );
  NAND2X1 U462 ( .A(\mem<11><4> ), .B(n985), .Y(n1624) );
  OAI21X1 U463 ( .A(n1033), .B(n985), .C(n1623), .Y(n1136) );
  NAND2X1 U464 ( .A(\mem<11><5> ), .B(n985), .Y(n1623) );
  OAI21X1 U465 ( .A(n1034), .B(n985), .C(n1622), .Y(n1135) );
  NAND2X1 U466 ( .A(\mem<11><6> ), .B(n985), .Y(n1622) );
  OAI21X1 U467 ( .A(n1035), .B(n985), .C(n1621), .Y(n1134) );
  NAND2X1 U468 ( .A(\mem<11><7> ), .B(n985), .Y(n1621) );
  NAND3X1 U469 ( .A(n973), .B(n1828), .C(n1620), .Y(n1629) );
  OAI21X1 U470 ( .A(n1036), .B(n984), .C(n1618), .Y(n1133) );
  NAND2X1 U471 ( .A(\mem<10><0> ), .B(n984), .Y(n1618) );
  OAI21X1 U472 ( .A(n1037), .B(n983), .C(n1617), .Y(n1132) );
  NAND2X1 U473 ( .A(\mem<10><1> ), .B(n984), .Y(n1617) );
  OAI21X1 U474 ( .A(n1038), .B(n983), .C(n1616), .Y(n1131) );
  NAND2X1 U475 ( .A(\mem<10><2> ), .B(n984), .Y(n1616) );
  OAI21X1 U476 ( .A(n1039), .B(n983), .C(n1615), .Y(n1130) );
  NAND2X1 U477 ( .A(\mem<10><3> ), .B(n984), .Y(n1615) );
  OAI21X1 U478 ( .A(n1040), .B(n983), .C(n1614), .Y(n1129) );
  NAND2X1 U479 ( .A(\mem<10><4> ), .B(n984), .Y(n1614) );
  OAI21X1 U480 ( .A(n1041), .B(n983), .C(n1613), .Y(n1128) );
  NAND2X1 U481 ( .A(\mem<10><5> ), .B(n984), .Y(n1613) );
  OAI21X1 U482 ( .A(n1042), .B(n983), .C(n1612), .Y(n1127) );
  NAND2X1 U483 ( .A(\mem<10><6> ), .B(n984), .Y(n1612) );
  OAI21X1 U484 ( .A(n1043), .B(n983), .C(n1611), .Y(n1126) );
  NAND2X1 U485 ( .A(\mem<10><7> ), .B(n984), .Y(n1611) );
  NAND3X1 U486 ( .A(n1766), .B(n1828), .C(n1651), .Y(n1619) );
  OAI21X1 U487 ( .A(n1028), .B(n982), .C(n1609), .Y(n1125) );
  NAND2X1 U488 ( .A(\mem<9><0> ), .B(n982), .Y(n1609) );
  OAI21X1 U489 ( .A(n1029), .B(n982), .C(n1608), .Y(n1124) );
  NAND2X1 U490 ( .A(\mem<9><1> ), .B(n982), .Y(n1608) );
  OAI21X1 U491 ( .A(n1030), .B(n982), .C(n1607), .Y(n1123) );
  NAND2X1 U492 ( .A(\mem<9><2> ), .B(n982), .Y(n1607) );
  OAI21X1 U493 ( .A(n1031), .B(n982), .C(n1606), .Y(n1122) );
  NAND2X1 U494 ( .A(\mem<9><3> ), .B(n982), .Y(n1606) );
  OAI21X1 U495 ( .A(n1032), .B(n982), .C(n1605), .Y(n1121) );
  NAND2X1 U496 ( .A(\mem<9><4> ), .B(n982), .Y(n1605) );
  OAI21X1 U497 ( .A(n1033), .B(n982), .C(n1604), .Y(n1120) );
  NAND2X1 U498 ( .A(\mem<9><5> ), .B(n982), .Y(n1604) );
  OAI21X1 U499 ( .A(n1034), .B(n982), .C(n1603), .Y(n1119) );
  NAND2X1 U500 ( .A(\mem<9><6> ), .B(n982), .Y(n1603) );
  OAI21X1 U501 ( .A(n1035), .B(n982), .C(n1602), .Y(n1118) );
  NAND2X1 U502 ( .A(\mem<9><7> ), .B(n982), .Y(n1602) );
  NAND3X1 U503 ( .A(n973), .B(n1828), .C(n1601), .Y(n1610) );
  OAI21X1 U504 ( .A(n1036), .B(n981), .C(n1599), .Y(n1117) );
  NAND2X1 U505 ( .A(\mem<8><0> ), .B(n981), .Y(n1599) );
  OAI21X1 U506 ( .A(n1037), .B(n980), .C(n1598), .Y(n1116) );
  NAND2X1 U507 ( .A(\mem<8><1> ), .B(n981), .Y(n1598) );
  OAI21X1 U508 ( .A(n1038), .B(n980), .C(n1597), .Y(n1115) );
  NAND2X1 U509 ( .A(\mem<8><2> ), .B(n981), .Y(n1597) );
  OAI21X1 U510 ( .A(n1039), .B(n980), .C(n1596), .Y(n1114) );
  NAND2X1 U511 ( .A(\mem<8><3> ), .B(n981), .Y(n1596) );
  OAI21X1 U512 ( .A(n1040), .B(n980), .C(n1595), .Y(n1113) );
  NAND2X1 U513 ( .A(\mem<8><4> ), .B(n981), .Y(n1595) );
  OAI21X1 U514 ( .A(n1041), .B(n980), .C(n1594), .Y(n1112) );
  NAND2X1 U515 ( .A(\mem<8><5> ), .B(n981), .Y(n1594) );
  OAI21X1 U516 ( .A(n1042), .B(n980), .C(n1593), .Y(n1111) );
  NAND2X1 U517 ( .A(\mem<8><6> ), .B(n981), .Y(n1593) );
  OAI21X1 U518 ( .A(n1043), .B(n980), .C(n1592), .Y(n1110) );
  NAND2X1 U519 ( .A(\mem<8><7> ), .B(n981), .Y(n1592) );
  NAND3X1 U520 ( .A(n1766), .B(n1828), .C(n1631), .Y(n1600) );
  OAI21X1 U521 ( .A(n1028), .B(n979), .C(n1589), .Y(n1109) );
  NAND2X1 U522 ( .A(\mem<7><0> ), .B(n979), .Y(n1589) );
  OAI21X1 U523 ( .A(n1029), .B(n979), .C(n1588), .Y(n1108) );
  NAND2X1 U524 ( .A(\mem<7><1> ), .B(n979), .Y(n1588) );
  OAI21X1 U525 ( .A(n1030), .B(n979), .C(n1587), .Y(n1107) );
  NAND2X1 U526 ( .A(\mem<7><2> ), .B(n979), .Y(n1587) );
  OAI21X1 U527 ( .A(n1031), .B(n979), .C(n1586), .Y(n1106) );
  NAND2X1 U528 ( .A(\mem<7><3> ), .B(n979), .Y(n1586) );
  OAI21X1 U529 ( .A(n1032), .B(n979), .C(n1585), .Y(n1105) );
  NAND2X1 U530 ( .A(\mem<7><4> ), .B(n979), .Y(n1585) );
  OAI21X1 U531 ( .A(n1033), .B(n979), .C(n1584), .Y(n1104) );
  NAND2X1 U532 ( .A(\mem<7><5> ), .B(n979), .Y(n1584) );
  OAI21X1 U533 ( .A(n1034), .B(n979), .C(n1583), .Y(n1103) );
  NAND2X1 U534 ( .A(\mem<7><6> ), .B(n979), .Y(n1583) );
  OAI21X1 U535 ( .A(n1035), .B(n979), .C(n1582), .Y(n1102) );
  NAND2X1 U536 ( .A(\mem<7><7> ), .B(n979), .Y(n1582) );
  NAND3X1 U537 ( .A(n973), .B(n1828), .C(n1581), .Y(n1590) );
  OAI21X1 U538 ( .A(n1036), .B(n978), .C(n1579), .Y(n1101) );
  NAND2X1 U539 ( .A(\mem<6><0> ), .B(n978), .Y(n1579) );
  OAI21X1 U540 ( .A(n1037), .B(n978), .C(n1578), .Y(n1100) );
  NAND2X1 U541 ( .A(\mem<6><1> ), .B(n978), .Y(n1578) );
  OAI21X1 U542 ( .A(n1038), .B(n978), .C(n1577), .Y(n1099) );
  NAND2X1 U543 ( .A(\mem<6><2> ), .B(n978), .Y(n1577) );
  OAI21X1 U544 ( .A(n1039), .B(n978), .C(n1576), .Y(n1098) );
  NAND2X1 U545 ( .A(\mem<6><3> ), .B(n978), .Y(n1576) );
  OAI21X1 U546 ( .A(n1040), .B(n978), .C(n1575), .Y(n1097) );
  NAND2X1 U547 ( .A(\mem<6><4> ), .B(n978), .Y(n1575) );
  OAI21X1 U548 ( .A(n1041), .B(n978), .C(n1574), .Y(n1096) );
  NAND2X1 U549 ( .A(\mem<6><5> ), .B(n978), .Y(n1574) );
  OAI21X1 U550 ( .A(n1042), .B(n978), .C(n1573), .Y(n1095) );
  NAND2X1 U551 ( .A(\mem<6><6> ), .B(n978), .Y(n1573) );
  OAI21X1 U552 ( .A(n1043), .B(n978), .C(n1572), .Y(n1094) );
  NAND2X1 U553 ( .A(\mem<6><7> ), .B(n978), .Y(n1572) );
  NAND3X1 U554 ( .A(n969), .B(n1828), .C(n1651), .Y(n1580) );
  OAI21X1 U555 ( .A(n1028), .B(n977), .C(n1570), .Y(n1093) );
  NAND2X1 U556 ( .A(\mem<5><0> ), .B(n977), .Y(n1570) );
  OAI21X1 U557 ( .A(n1029), .B(n977), .C(n1569), .Y(n1092) );
  NAND2X1 U558 ( .A(\mem<5><1> ), .B(n977), .Y(n1569) );
  OAI21X1 U559 ( .A(n1030), .B(n977), .C(n1568), .Y(n1091) );
  NAND2X1 U560 ( .A(\mem<5><2> ), .B(n977), .Y(n1568) );
  OAI21X1 U561 ( .A(n1031), .B(n977), .C(n1567), .Y(n1090) );
  NAND2X1 U562 ( .A(\mem<5><3> ), .B(n977), .Y(n1567) );
  OAI21X1 U563 ( .A(n1032), .B(n977), .C(n1566), .Y(n1089) );
  NAND2X1 U564 ( .A(\mem<5><4> ), .B(n977), .Y(n1566) );
  OAI21X1 U565 ( .A(n1033), .B(n977), .C(n1565), .Y(n1088) );
  NAND2X1 U566 ( .A(\mem<5><5> ), .B(n977), .Y(n1565) );
  OAI21X1 U567 ( .A(n1034), .B(n977), .C(n1564), .Y(n1087) );
  NAND2X1 U568 ( .A(\mem<5><6> ), .B(n977), .Y(n1564) );
  OAI21X1 U569 ( .A(n1035), .B(n977), .C(n1563), .Y(n1086) );
  NAND2X1 U570 ( .A(\mem<5><7> ), .B(n977), .Y(n1563) );
  NAND3X1 U571 ( .A(n973), .B(n1828), .C(n1562), .Y(n1571) );
  OAI21X1 U572 ( .A(n1036), .B(n976), .C(n1560), .Y(n1085) );
  NAND2X1 U573 ( .A(\mem<4><0> ), .B(n976), .Y(n1560) );
  OAI21X1 U574 ( .A(n1037), .B(n976), .C(n1559), .Y(n1084) );
  NAND2X1 U575 ( .A(\mem<4><1> ), .B(n976), .Y(n1559) );
  OAI21X1 U576 ( .A(n1038), .B(n976), .C(n1558), .Y(n1083) );
  NAND2X1 U577 ( .A(\mem<4><2> ), .B(n976), .Y(n1558) );
  OAI21X1 U578 ( .A(n1039), .B(n976), .C(n1557), .Y(n1082) );
  NAND2X1 U579 ( .A(\mem<4><3> ), .B(n976), .Y(n1557) );
  OAI21X1 U580 ( .A(n1040), .B(n976), .C(n1556), .Y(n1081) );
  NAND2X1 U581 ( .A(\mem<4><4> ), .B(n976), .Y(n1556) );
  OAI21X1 U582 ( .A(n1041), .B(n976), .C(n1555), .Y(n1080) );
  NAND2X1 U583 ( .A(\mem<4><5> ), .B(n976), .Y(n1555) );
  OAI21X1 U584 ( .A(n1042), .B(n976), .C(n1554), .Y(n1079) );
  NAND2X1 U585 ( .A(\mem<4><6> ), .B(n976), .Y(n1554) );
  OAI21X1 U586 ( .A(n1043), .B(n976), .C(n1553), .Y(n1078) );
  NAND2X1 U587 ( .A(\mem<4><7> ), .B(n976), .Y(n1553) );
  NAND3X1 U588 ( .A(n969), .B(n1828), .C(n1631), .Y(n1561) );
  OAI21X1 U590 ( .A(n1028), .B(n975), .C(n1550), .Y(n1077) );
  NAND2X1 U591 ( .A(\mem<3><0> ), .B(n975), .Y(n1550) );
  OAI21X1 U592 ( .A(n1029), .B(n975), .C(n1549), .Y(n1076) );
  NAND2X1 U593 ( .A(\mem<3><1> ), .B(n975), .Y(n1549) );
  OAI21X1 U594 ( .A(n1030), .B(n975), .C(n1548), .Y(n1075) );
  NAND2X1 U595 ( .A(\mem<3><2> ), .B(n975), .Y(n1548) );
  OAI21X1 U596 ( .A(n1031), .B(n975), .C(n1547), .Y(n1074) );
  NAND2X1 U597 ( .A(\mem<3><3> ), .B(n975), .Y(n1547) );
  OAI21X1 U598 ( .A(n1032), .B(n975), .C(n1546), .Y(n1073) );
  NAND2X1 U599 ( .A(\mem<3><4> ), .B(n975), .Y(n1546) );
  OAI21X1 U600 ( .A(n1033), .B(n975), .C(n1545), .Y(n1072) );
  NAND2X1 U601 ( .A(\mem<3><5> ), .B(n975), .Y(n1545) );
  OAI21X1 U602 ( .A(n1034), .B(n975), .C(n1544), .Y(n1071) );
  NAND2X1 U603 ( .A(\mem<3><6> ), .B(n975), .Y(n1544) );
  OAI21X1 U604 ( .A(n1035), .B(n975), .C(n1543), .Y(n1070) );
  NAND2X1 U605 ( .A(\mem<3><7> ), .B(n975), .Y(n1543) );
  NAND3X1 U606 ( .A(n973), .B(n1828), .C(n1542), .Y(n1551) );
  OAI21X1 U607 ( .A(n1036), .B(n974), .C(n1540), .Y(n1069) );
  NAND2X1 U608 ( .A(\mem<2><0> ), .B(n974), .Y(n1540) );
  OAI21X1 U609 ( .A(n1037), .B(n974), .C(n1539), .Y(n1068) );
  NAND2X1 U610 ( .A(\mem<2><1> ), .B(n974), .Y(n1539) );
  OAI21X1 U611 ( .A(n1038), .B(n974), .C(n1538), .Y(n1067) );
  NAND2X1 U612 ( .A(\mem<2><2> ), .B(n974), .Y(n1538) );
  OAI21X1 U613 ( .A(n1039), .B(n974), .C(n1537), .Y(n1066) );
  NAND2X1 U614 ( .A(\mem<2><3> ), .B(n974), .Y(n1537) );
  OAI21X1 U615 ( .A(n1040), .B(n974), .C(n1536), .Y(n1065) );
  NAND2X1 U616 ( .A(\mem<2><4> ), .B(n974), .Y(n1536) );
  OAI21X1 U617 ( .A(n1041), .B(n974), .C(n1535), .Y(n1064) );
  NAND2X1 U618 ( .A(\mem<2><5> ), .B(n974), .Y(n1535) );
  OAI21X1 U619 ( .A(n1042), .B(n974), .C(n1534), .Y(n1063) );
  NAND2X1 U620 ( .A(\mem<2><6> ), .B(n974), .Y(n1534) );
  OAI21X1 U621 ( .A(n1043), .B(n974), .C(n1533), .Y(n1062) );
  NAND2X1 U622 ( .A(\mem<2><7> ), .B(n974), .Y(n1533) );
  NAND3X1 U623 ( .A(n967), .B(n1828), .C(n1651), .Y(n1541) );
  OAI21X1 U624 ( .A(n1028), .B(n8), .C(n1532), .Y(n1061) );
  NAND2X1 U625 ( .A(\mem<1><0> ), .B(n8), .Y(n1532) );
  OAI21X1 U626 ( .A(n1029), .B(n8), .C(n1531), .Y(n1060) );
  NAND2X1 U627 ( .A(\mem<1><1> ), .B(n8), .Y(n1531) );
  OAI21X1 U628 ( .A(n1030), .B(n8), .C(n1530), .Y(n1059) );
  NAND2X1 U629 ( .A(\mem<1><2> ), .B(n8), .Y(n1530) );
  OAI21X1 U630 ( .A(n1031), .B(n8), .C(n1529), .Y(n1058) );
  NAND2X1 U631 ( .A(\mem<1><3> ), .B(n8), .Y(n1529) );
  OAI21X1 U632 ( .A(n1032), .B(n8), .C(n1528), .Y(n1057) );
  NAND2X1 U633 ( .A(\mem<1><4> ), .B(n8), .Y(n1528) );
  OAI21X1 U634 ( .A(n1033), .B(n8), .C(n1527), .Y(n1056) );
  NAND2X1 U635 ( .A(\mem<1><5> ), .B(n8), .Y(n1527) );
  OAI21X1 U636 ( .A(n1034), .B(n8), .C(n1526), .Y(n1055) );
  NAND2X1 U637 ( .A(\mem<1><6> ), .B(n8), .Y(n1526) );
  OAI21X1 U638 ( .A(n1035), .B(n8), .C(n1525), .Y(n1054) );
  NAND2X1 U639 ( .A(\mem<1><7> ), .B(n8), .Y(n1525) );
  NOR2X1 U641 ( .A(n965), .B(\addr_1c<4> ), .Y(n1818) );
  OAI21X1 U642 ( .A(n1036), .B(n972), .C(n1522), .Y(n1053) );
  NAND2X1 U643 ( .A(\mem<0><0> ), .B(n972), .Y(n1522) );
  OAI21X1 U644 ( .A(n1037), .B(n972), .C(n1521), .Y(n1052) );
  NAND2X1 U645 ( .A(\mem<0><1> ), .B(n972), .Y(n1521) );
  OAI21X1 U646 ( .A(n1038), .B(n972), .C(n1520), .Y(n1051) );
  NAND2X1 U647 ( .A(\mem<0><2> ), .B(n972), .Y(n1520) );
  OAI21X1 U648 ( .A(n1039), .B(n972), .C(n1519), .Y(n1050) );
  NAND2X1 U649 ( .A(\mem<0><3> ), .B(n972), .Y(n1519) );
  OAI21X1 U650 ( .A(n1040), .B(n972), .C(n1518), .Y(n1049) );
  NAND2X1 U651 ( .A(\mem<0><4> ), .B(n972), .Y(n1518) );
  OAI21X1 U652 ( .A(n1041), .B(n972), .C(n1517), .Y(n1048) );
  NAND2X1 U653 ( .A(\mem<0><5> ), .B(n972), .Y(n1517) );
  OAI21X1 U654 ( .A(n1042), .B(n972), .C(n1516), .Y(n1047) );
  NAND2X1 U655 ( .A(\mem<0><6> ), .B(n972), .Y(n1516) );
  OAI21X1 U656 ( .A(n1043), .B(n972), .C(n1515), .Y(n1046) );
  NAND2X1 U657 ( .A(\mem<0><7> ), .B(n972), .Y(n1515) );
  NAND3X1 U658 ( .A(n967), .B(n1828), .C(n1631), .Y(n1523) );
  NOR3X1 U661 ( .A(n1511), .B(\addr_1c<7> ), .C(\addr_1c<6> ), .Y(n1512) );
  NOR3X1 U662 ( .A(n1510), .B(\addr_1c<11> ), .C(\addr_1c<10> ), .Y(n1513) );
  AOI21X1 U663 ( .A(n461), .B(n1509), .C(n963), .Y(n1838) );
  OAI21X1 U665 ( .A(rd), .B(n1508), .C(wr), .Y(n1509) );
  NAND3X1 U667 ( .A(n1507), .B(n1023), .C(n1506), .Y(n1508) );
  NOR3X1 U668 ( .A(rd1), .B(rd3), .C(rd2), .Y(n1506) );
  NOR2X1 U669 ( .A(wr3), .B(wr2), .Y(n1507) );
  AOI21X1 U670 ( .A(n448), .B(n1504), .C(n1014), .Y(\data_out_1c<9> ) );
  NOR3X1 U671 ( .A(n2), .B(n1503), .C(n4), .Y(n1504) );
  AOI22X1 U673 ( .A(\mem<16><1> ), .B(n1786), .C(\mem<0><1> ), .D(n1631), .Y(
        n1501) );
  AOI22X1 U674 ( .A(\mem<18><1> ), .B(n1806), .C(\mem<2><1> ), .D(n1651), .Y(
        n1502) );
  AOI22X1 U676 ( .A(\mem<20><1> ), .B(n1786), .C(\mem<4><1> ), .D(n1631), .Y(
        n1499) );
  AOI22X1 U677 ( .A(\mem<22><1> ), .B(n1806), .C(\mem<6><1> ), .D(n1651), .Y(
        n1500) );
  AOI22X1 U678 ( .A(n1591), .B(n892), .C(n1630), .D(n932), .Y(n1505) );
  AOI22X1 U680 ( .A(\mem<28><1> ), .B(n1786), .C(\mem<12><1> ), .D(n1631), .Y(
        n1497) );
  AOI22X1 U681 ( .A(\mem<30><1> ), .B(n1806), .C(\mem<14><1> ), .D(n1651), .Y(
        n1498) );
  AOI22X1 U683 ( .A(\mem<24><1> ), .B(n1786), .C(\mem<8><1> ), .D(n1631), .Y(
        n1495) );
  AOI22X1 U684 ( .A(\mem<26><1> ), .B(n1806), .C(\mem<10><1> ), .D(n1651), .Y(
        n1496) );
  AOI21X1 U685 ( .A(n447), .B(n1493), .C(n1014), .Y(\data_out_1c<8> ) );
  NOR3X1 U686 ( .A(n939), .B(n1491), .C(n950), .Y(n1493) );
  AOI21X1 U687 ( .A(n1489), .B(n1488), .C(n971), .Y(n1490) );
  AOI22X1 U688 ( .A(\mem<16><0> ), .B(n1786), .C(\mem<0><0> ), .D(n1631), .Y(
        n1488) );
  AOI22X1 U689 ( .A(\mem<18><0> ), .B(n1806), .C(\mem<2><0> ), .D(n1651), .Y(
        n1489) );
  AOI21X1 U690 ( .A(n1487), .B(n1486), .C(n970), .Y(n1492) );
  AOI22X1 U691 ( .A(\mem<20><0> ), .B(n1786), .C(\mem<4><0> ), .D(n1631), .Y(
        n1486) );
  AOI22X1 U692 ( .A(\mem<22><0> ), .B(n1806), .C(\mem<6><0> ), .D(n1651), .Y(
        n1487) );
  AOI22X1 U693 ( .A(n1591), .B(n890), .C(n1630), .D(n930), .Y(n1494) );
  AOI22X1 U695 ( .A(\mem<28><0> ), .B(n1786), .C(\mem<12><0> ), .D(n1631), .Y(
        n1484) );
  AOI22X1 U696 ( .A(\mem<30><0> ), .B(n1806), .C(\mem<14><0> ), .D(n1651), .Y(
        n1485) );
  AOI22X1 U698 ( .A(\mem<24><0> ), .B(n1786), .C(\mem<8><0> ), .D(n1631), .Y(
        n1482) );
  AOI22X1 U699 ( .A(\mem<26><0> ), .B(n1806), .C(\mem<10><0> ), .D(n1651), .Y(
        n1483) );
  OAI21X1 U700 ( .A(n23), .B(n50), .C(rd1), .Y(n1481) );
  AOI22X1 U702 ( .A(\mem<17><7> ), .B(n1680), .C(\mem<19><7> ), .D(n1699), .Y(
        n1476) );
  AOI22X1 U703 ( .A(\mem<21><7> ), .B(n1718), .C(\mem<23><7> ), .D(n1737), .Y(
        n1477) );
  AOI22X1 U704 ( .A(\mem<25><7> ), .B(n1756), .C(\mem<27><7> ), .D(n1776), .Y(
        n1479) );
  AOI22X1 U705 ( .A(\mem<29><7> ), .B(n1796), .C(\mem<31><7> ), .D(n1817), .Y(
        n1480) );
  AOI22X1 U707 ( .A(\mem<1><7> ), .B(n1524), .C(\mem<3><7> ), .D(n1542), .Y(
        n1471) );
  AOI22X1 U708 ( .A(\mem<5><7> ), .B(n1562), .C(\mem<7><7> ), .D(n1581), .Y(
        n1472) );
  AOI22X1 U709 ( .A(\mem<9><7> ), .B(n1601), .C(\mem<11><7> ), .D(n1620), .Y(
        n1474) );
  AOI22X1 U710 ( .A(\mem<13><7> ), .B(n1641), .C(\mem<15><7> ), .D(n1661), .Y(
        n1475) );
  OAI21X1 U711 ( .A(n21), .B(n37), .C(rd1), .Y(n1470) );
  AOI22X1 U713 ( .A(\mem<17><6> ), .B(n1680), .C(\mem<19><6> ), .D(n1699), .Y(
        n1465) );
  AOI22X1 U714 ( .A(\mem<21><6> ), .B(n1718), .C(\mem<23><6> ), .D(n1737), .Y(
        n1466) );
  AOI22X1 U715 ( .A(\mem<25><6> ), .B(n1756), .C(\mem<27><6> ), .D(n1776), .Y(
        n1468) );
  AOI22X1 U716 ( .A(\mem<29><6> ), .B(n1796), .C(\mem<31><6> ), .D(n1817), .Y(
        n1469) );
  AOI22X1 U718 ( .A(\mem<1><6> ), .B(n1524), .C(\mem<3><6> ), .D(n1542), .Y(
        n1460) );
  AOI22X1 U719 ( .A(\mem<5><6> ), .B(n1562), .C(\mem<7><6> ), .D(n1581), .Y(
        n1461) );
  AOI22X1 U720 ( .A(\mem<9><6> ), .B(n1601), .C(\mem<11><6> ), .D(n1620), .Y(
        n1463) );
  AOI22X1 U721 ( .A(\mem<13><6> ), .B(n1641), .C(\mem<15><6> ), .D(n1661), .Y(
        n1464) );
  OAI21X1 U722 ( .A(n19), .B(n35), .C(rd1), .Y(n1459) );
  AOI22X1 U724 ( .A(\mem<17><5> ), .B(n1680), .C(\mem<19><5> ), .D(n1699), .Y(
        n1454) );
  AOI22X1 U725 ( .A(\mem<21><5> ), .B(n1718), .C(\mem<23><5> ), .D(n1737), .Y(
        n1455) );
  AOI22X1 U726 ( .A(\mem<25><5> ), .B(n1756), .C(\mem<27><5> ), .D(n1776), .Y(
        n1457) );
  AOI22X1 U727 ( .A(\mem<29><5> ), .B(n1796), .C(\mem<31><5> ), .D(n1817), .Y(
        n1458) );
  AOI22X1 U729 ( .A(\mem<1><5> ), .B(n1524), .C(\mem<3><5> ), .D(n1542), .Y(
        n1449) );
  AOI22X1 U730 ( .A(\mem<5><5> ), .B(n1562), .C(\mem<7><5> ), .D(n1581), .Y(
        n1450) );
  AOI22X1 U731 ( .A(\mem<9><5> ), .B(n1601), .C(\mem<11><5> ), .D(n1620), .Y(
        n1452) );
  AOI22X1 U732 ( .A(\mem<13><5> ), .B(n1641), .C(\mem<15><5> ), .D(n1661), .Y(
        n1453) );
  OAI21X1 U733 ( .A(n17), .B(n33), .C(rd1), .Y(n1448) );
  AOI22X1 U735 ( .A(\mem<17><4> ), .B(n1680), .C(\mem<19><4> ), .D(n1699), .Y(
        n1443) );
  AOI22X1 U736 ( .A(\mem<21><4> ), .B(n1718), .C(\mem<23><4> ), .D(n1737), .Y(
        n1444) );
  AOI22X1 U737 ( .A(\mem<25><4> ), .B(n1756), .C(\mem<27><4> ), .D(n1776), .Y(
        n1446) );
  AOI22X1 U738 ( .A(\mem<29><4> ), .B(n1796), .C(\mem<31><4> ), .D(n1817), .Y(
        n1447) );
  AOI22X1 U740 ( .A(\mem<1><4> ), .B(n1524), .C(\mem<3><4> ), .D(n1542), .Y(
        n1438) );
  AOI22X1 U741 ( .A(\mem<5><4> ), .B(n1562), .C(\mem<7><4> ), .D(n1581), .Y(
        n1439) );
  AOI22X1 U742 ( .A(\mem<9><4> ), .B(n1601), .C(\mem<11><4> ), .D(n1620), .Y(
        n1441) );
  AOI22X1 U743 ( .A(\mem<13><4> ), .B(n1641), .C(\mem<15><4> ), .D(n1661), .Y(
        n1442) );
  OAI21X1 U744 ( .A(n15), .B(n31), .C(rd1), .Y(n1437) );
  AOI22X1 U746 ( .A(\mem<17><3> ), .B(n1680), .C(\mem<19><3> ), .D(n1699), .Y(
        n1432) );
  AOI22X1 U747 ( .A(\mem<21><3> ), .B(n1718), .C(\mem<23><3> ), .D(n1737), .Y(
        n1433) );
  AOI22X1 U748 ( .A(\mem<25><3> ), .B(n1756), .C(\mem<27><3> ), .D(n1776), .Y(
        n1435) );
  AOI22X1 U749 ( .A(\mem<29><3> ), .B(n1796), .C(\mem<31><3> ), .D(n1817), .Y(
        n1436) );
  AOI22X1 U751 ( .A(\mem<1><3> ), .B(n1524), .C(\mem<3><3> ), .D(n1542), .Y(
        n1427) );
  AOI22X1 U752 ( .A(\mem<5><3> ), .B(n1562), .C(\mem<7><3> ), .D(n1581), .Y(
        n1428) );
  AOI22X1 U753 ( .A(\mem<9><3> ), .B(n1601), .C(\mem<11><3> ), .D(n1620), .Y(
        n1430) );
  AOI22X1 U754 ( .A(\mem<13><3> ), .B(n1641), .C(\mem<15><3> ), .D(n1661), .Y(
        n1431) );
  OAI21X1 U755 ( .A(n13), .B(n29), .C(rd1), .Y(n1426) );
  AOI22X1 U757 ( .A(\mem<17><2> ), .B(n1680), .C(\mem<19><2> ), .D(n1699), .Y(
        n1421) );
  AOI22X1 U758 ( .A(\mem<21><2> ), .B(n1718), .C(\mem<23><2> ), .D(n1737), .Y(
        n1422) );
  AOI22X1 U759 ( .A(\mem<25><2> ), .B(n1756), .C(\mem<27><2> ), .D(n1776), .Y(
        n1424) );
  AOI22X1 U760 ( .A(\mem<29><2> ), .B(n1796), .C(\mem<31><2> ), .D(n1817), .Y(
        n1425) );
  AOI22X1 U762 ( .A(\mem<1><2> ), .B(n1524), .C(\mem<3><2> ), .D(n1542), .Y(
        n1416) );
  AOI22X1 U763 ( .A(\mem<5><2> ), .B(n1562), .C(\mem<7><2> ), .D(n1581), .Y(
        n1417) );
  AOI22X1 U764 ( .A(\mem<9><2> ), .B(n1601), .C(\mem<11><2> ), .D(n1620), .Y(
        n1419) );
  AOI22X1 U765 ( .A(\mem<13><2> ), .B(n1641), .C(\mem<15><2> ), .D(n1661), .Y(
        n1420) );
  OAI21X1 U766 ( .A(n11), .B(n27), .C(rd1), .Y(n1415) );
  AOI22X1 U768 ( .A(\mem<17><1> ), .B(n1680), .C(\mem<19><1> ), .D(n1699), .Y(
        n1410) );
  AOI22X1 U769 ( .A(\mem<21><1> ), .B(n1718), .C(\mem<23><1> ), .D(n1737), .Y(
        n1411) );
  AOI22X1 U770 ( .A(\mem<25><1> ), .B(n1756), .C(\mem<27><1> ), .D(n1776), .Y(
        n1413) );
  AOI22X1 U771 ( .A(\mem<29><1> ), .B(n1796), .C(\mem<31><1> ), .D(n1817), .Y(
        n1414) );
  AOI22X1 U773 ( .A(\mem<1><1> ), .B(n1524), .C(\mem<3><1> ), .D(n1542), .Y(
        n1405) );
  AOI22X1 U774 ( .A(\mem<5><1> ), .B(n1562), .C(\mem<7><1> ), .D(n1581), .Y(
        n1406) );
  AOI22X1 U775 ( .A(\mem<9><1> ), .B(n1601), .C(\mem<11><1> ), .D(n1620), .Y(
        n1408) );
  AOI22X1 U776 ( .A(\mem<13><1> ), .B(n1641), .C(\mem<15><1> ), .D(n1661), .Y(
        n1409) );
  AOI21X1 U777 ( .A(n435), .B(n1403), .C(n1014), .Y(\data_out_1c<15> ) );
  NOR3X1 U778 ( .A(n938), .B(n1401), .C(n949), .Y(n1403) );
  AOI21X1 U779 ( .A(n1399), .B(n1398), .C(n971), .Y(n1400) );
  AOI22X1 U780 ( .A(\mem<16><7> ), .B(n1786), .C(\mem<0><7> ), .D(n1631), .Y(
        n1398) );
  AOI22X1 U781 ( .A(\mem<18><7> ), .B(n1806), .C(\mem<2><7> ), .D(n1651), .Y(
        n1399) );
  AOI21X1 U782 ( .A(n1397), .B(n1396), .C(n970), .Y(n1402) );
  AOI22X1 U783 ( .A(\mem<20><7> ), .B(n1786), .C(\mem<4><7> ), .D(n1631), .Y(
        n1396) );
  AOI22X1 U784 ( .A(\mem<22><7> ), .B(n1806), .C(\mem<6><7> ), .D(n1651), .Y(
        n1397) );
  AOI22X1 U785 ( .A(n1591), .B(n888), .C(n1630), .D(n928), .Y(n1404) );
  AOI22X1 U787 ( .A(\mem<28><7> ), .B(n1786), .C(\mem<12><7> ), .D(n1631), .Y(
        n1394) );
  AOI22X1 U788 ( .A(\mem<30><7> ), .B(n1806), .C(\mem<14><7> ), .D(n1651), .Y(
        n1395) );
  AOI22X1 U790 ( .A(\mem<24><7> ), .B(n1786), .C(\mem<8><7> ), .D(n1631), .Y(
        n1392) );
  AOI22X1 U791 ( .A(\mem<26><7> ), .B(n1806), .C(\mem<10><7> ), .D(n1651), .Y(
        n1393) );
  AOI21X1 U792 ( .A(n434), .B(n1390), .C(n1014), .Y(\data_out_1c<14> ) );
  NOR3X1 U793 ( .A(n937), .B(n1388), .C(n948), .Y(n1390) );
  AOI21X1 U794 ( .A(n1386), .B(n1385), .C(n971), .Y(n1387) );
  AOI22X1 U795 ( .A(\mem<16><6> ), .B(n1786), .C(\mem<0><6> ), .D(n1631), .Y(
        n1385) );
  AOI22X1 U796 ( .A(\mem<18><6> ), .B(n1806), .C(\mem<2><6> ), .D(n1651), .Y(
        n1386) );
  AOI21X1 U797 ( .A(n1384), .B(n1383), .C(n970), .Y(n1389) );
  AOI22X1 U798 ( .A(\mem<20><6> ), .B(n1786), .C(\mem<4><6> ), .D(n1631), .Y(
        n1383) );
  AOI22X1 U799 ( .A(\mem<22><6> ), .B(n1806), .C(\mem<6><6> ), .D(n1651), .Y(
        n1384) );
  AOI22X1 U800 ( .A(n1591), .B(n886), .C(n1630), .D(n926), .Y(n1391) );
  AOI22X1 U802 ( .A(\mem<28><6> ), .B(n1786), .C(\mem<12><6> ), .D(n1631), .Y(
        n1381) );
  AOI22X1 U803 ( .A(\mem<30><6> ), .B(n1806), .C(\mem<14><6> ), .D(n1651), .Y(
        n1382) );
  AOI22X1 U805 ( .A(\mem<24><6> ), .B(n1786), .C(\mem<8><6> ), .D(n1631), .Y(
        n1379) );
  AOI22X1 U806 ( .A(\mem<26><6> ), .B(n1806), .C(\mem<10><6> ), .D(n1651), .Y(
        n1380) );
  AOI21X1 U807 ( .A(n422), .B(n1377), .C(n1014), .Y(\data_out_1c<13> ) );
  NOR3X1 U808 ( .A(n936), .B(n1375), .C(n947), .Y(n1377) );
  AOI21X1 U809 ( .A(n1373), .B(n1372), .C(n971), .Y(n1374) );
  AOI22X1 U810 ( .A(\mem<16><5> ), .B(n1786), .C(\mem<0><5> ), .D(n1631), .Y(
        n1372) );
  AOI22X1 U811 ( .A(\mem<18><5> ), .B(n1806), .C(\mem<2><5> ), .D(n1651), .Y(
        n1373) );
  AOI21X1 U812 ( .A(n1371), .B(n1370), .C(n970), .Y(n1376) );
  AOI22X1 U813 ( .A(\mem<20><5> ), .B(n1786), .C(\mem<4><5> ), .D(n1631), .Y(
        n1370) );
  AOI22X1 U814 ( .A(\mem<22><5> ), .B(n1806), .C(\mem<6><5> ), .D(n1651), .Y(
        n1371) );
  AOI22X1 U815 ( .A(n1591), .B(n884), .C(n1630), .D(n924), .Y(n1378) );
  AOI22X1 U817 ( .A(\mem<28><5> ), .B(n1786), .C(\mem<12><5> ), .D(n1631), .Y(
        n1368) );
  AOI22X1 U818 ( .A(\mem<30><5> ), .B(n1806), .C(\mem<14><5> ), .D(n1651), .Y(
        n1369) );
  AOI22X1 U820 ( .A(\mem<24><5> ), .B(n1786), .C(\mem<8><5> ), .D(n1631), .Y(
        n1366) );
  AOI22X1 U821 ( .A(\mem<26><5> ), .B(n1806), .C(\mem<10><5> ), .D(n1651), .Y(
        n1367) );
  AOI21X1 U822 ( .A(n421), .B(n1364), .C(n1014), .Y(\data_out_1c<12> ) );
  NOR3X1 U823 ( .A(n935), .B(n1362), .C(n946), .Y(n1364) );
  AOI21X1 U824 ( .A(n1360), .B(n1359), .C(n971), .Y(n1361) );
  AOI22X1 U825 ( .A(\mem<16><4> ), .B(n1786), .C(\mem<0><4> ), .D(n1631), .Y(
        n1359) );
  AOI22X1 U826 ( .A(\mem<18><4> ), .B(n1806), .C(\mem<2><4> ), .D(n1651), .Y(
        n1360) );
  AOI21X1 U827 ( .A(n1358), .B(n1357), .C(n970), .Y(n1363) );
  AOI22X1 U828 ( .A(\mem<20><4> ), .B(n1786), .C(\mem<4><4> ), .D(n1631), .Y(
        n1357) );
  AOI22X1 U829 ( .A(\mem<22><4> ), .B(n1806), .C(\mem<6><4> ), .D(n1651), .Y(
        n1358) );
  AOI22X1 U830 ( .A(n1591), .B(n882), .C(n1630), .D(n922), .Y(n1365) );
  AOI22X1 U832 ( .A(\mem<28><4> ), .B(n1786), .C(\mem<12><4> ), .D(n1631), .Y(
        n1355) );
  AOI22X1 U833 ( .A(\mem<30><4> ), .B(n1806), .C(\mem<14><4> ), .D(n1651), .Y(
        n1356) );
  AOI22X1 U835 ( .A(\mem<24><4> ), .B(n1786), .C(\mem<8><4> ), .D(n1631), .Y(
        n1353) );
  AOI22X1 U836 ( .A(\mem<26><4> ), .B(n1806), .C(\mem<10><4> ), .D(n1651), .Y(
        n1354) );
  AOI21X1 U837 ( .A(n409), .B(n1351), .C(n1014), .Y(\data_out_1c<11> ) );
  NOR3X1 U838 ( .A(n934), .B(n1349), .C(n945), .Y(n1351) );
  AOI21X1 U839 ( .A(n1347), .B(n1346), .C(n971), .Y(n1348) );
  AOI22X1 U840 ( .A(\mem<16><3> ), .B(n1786), .C(\mem<0><3> ), .D(n1631), .Y(
        n1346) );
  AOI22X1 U841 ( .A(\mem<18><3> ), .B(n1806), .C(\mem<2><3> ), .D(n1651), .Y(
        n1347) );
  AOI21X1 U842 ( .A(n1345), .B(n1344), .C(n970), .Y(n1350) );
  AOI22X1 U843 ( .A(\mem<20><3> ), .B(n1786), .C(\mem<4><3> ), .D(n1631), .Y(
        n1344) );
  AOI22X1 U844 ( .A(\mem<22><3> ), .B(n1806), .C(\mem<6><3> ), .D(n1651), .Y(
        n1345) );
  AOI22X1 U845 ( .A(n1591), .B(n880), .C(n1630), .D(n920), .Y(n1352) );
  AOI22X1 U847 ( .A(\mem<28><3> ), .B(n1786), .C(\mem<12><3> ), .D(n1631), .Y(
        n1342) );
  AOI22X1 U848 ( .A(\mem<30><3> ), .B(n1806), .C(\mem<14><3> ), .D(n1651), .Y(
        n1343) );
  AOI22X1 U850 ( .A(\mem<24><3> ), .B(n1786), .C(\mem<8><3> ), .D(n1631), .Y(
        n1340) );
  AOI22X1 U851 ( .A(\mem<26><3> ), .B(n1806), .C(\mem<10><3> ), .D(n1651), .Y(
        n1341) );
  AOI21X1 U852 ( .A(n408), .B(n1338), .C(n1014), .Y(\data_out_1c<10> ) );
  NOR3X1 U853 ( .A(n933), .B(n1336), .C(n944), .Y(n1338) );
  AOI21X1 U854 ( .A(n1334), .B(n1333), .C(n971), .Y(n1335) );
  AOI22X1 U855 ( .A(\mem<16><2> ), .B(n1786), .C(\mem<0><2> ), .D(n1631), .Y(
        n1333) );
  AOI22X1 U856 ( .A(\mem<18><2> ), .B(n1806), .C(\mem<2><2> ), .D(n1651), .Y(
        n1334) );
  AOI21X1 U857 ( .A(n1332), .B(n1331), .C(n970), .Y(n1337) );
  AOI22X1 U858 ( .A(\mem<20><2> ), .B(n1786), .C(\mem<4><2> ), .D(n1631), .Y(
        n1331) );
  AOI22X1 U859 ( .A(\mem<22><2> ), .B(n1806), .C(\mem<6><2> ), .D(n1651), .Y(
        n1332) );
  AOI22X1 U860 ( .A(n1591), .B(n878), .C(n1630), .D(n918), .Y(n1339) );
  AOI22X1 U862 ( .A(\mem<28><2> ), .B(n1786), .C(\mem<12><2> ), .D(n1631), .Y(
        n1329) );
  AOI22X1 U863 ( .A(\mem<30><2> ), .B(n1806), .C(\mem<14><2> ), .D(n1651), .Y(
        n1330) );
  AOI22X1 U865 ( .A(\mem<24><2> ), .B(n1786), .C(\mem<8><2> ), .D(n1631), .Y(
        n1327) );
  AOI22X1 U866 ( .A(\mem<26><2> ), .B(n1806), .C(\mem<10><2> ), .D(n1651), .Y(
        n1328) );
  NOR2X1 U867 ( .A(\addr_1c<3> ), .B(\addr_1c<4> ), .Y(n1326) );
  NOR2X1 U868 ( .A(n1027), .B(\addr_1c<4> ), .Y(n1325) );
  OAI21X1 U869 ( .A(n9), .B(n25), .C(rd1), .Y(n1324) );
  AOI22X1 U871 ( .A(\mem<17><0> ), .B(n1680), .C(\mem<19><0> ), .D(n1699), .Y(
        n1319) );
  AOI22X1 U872 ( .A(\mem<21><0> ), .B(n1718), .C(\mem<23><0> ), .D(n1737), .Y(
        n1320) );
  AOI22X1 U873 ( .A(\mem<25><0> ), .B(n1756), .C(\mem<27><0> ), .D(n1776), .Y(
        n1322) );
  AOI22X1 U874 ( .A(\mem<29><0> ), .B(n1796), .C(\mem<31><0> ), .D(n1817), .Y(
        n1323) );
  AOI22X1 U876 ( .A(\mem<1><0> ), .B(n1524), .C(\mem<3><0> ), .D(n1542), .Y(
        n1312) );
  NAND2X1 U877 ( .A(n1025), .B(n1026), .Y(n1514) );
  AOI22X1 U878 ( .A(\mem<5><0> ), .B(n1562), .C(\mem<7><0> ), .D(n1581), .Y(
        n1313) );
  NAND2X1 U879 ( .A(\addr_1c<1> ), .B(n1026), .Y(n1552) );
  AOI22X1 U880 ( .A(\mem<9><0> ), .B(n1601), .C(\mem<11><0> ), .D(n1620), .Y(
        n1315) );
  AOI22X1 U881 ( .A(\mem<13><0> ), .B(n1641), .C(\mem<15><0> ), .D(n1661), .Y(
        n1316) );
  dff_156 ff0 ( .q(rd1), .d(rd0), .clk(clk), .rst(n1012) );
  dff_155 ff1 ( .q(wr1), .d(wr0), .clk(clk), .rst(n1012) );
  dff_154 \reg0[0]  ( .q(\addr_1c<0> ), .d(\addr<0> ), .clk(clk), .rst(n1012)
         );
  dff_153 \reg0[1]  ( .q(\addr_1c<1> ), .d(\addr<1> ), .clk(clk), .rst(n1012)
         );
  dff_152 \reg0[2]  ( .q(\addr_1c<2> ), .d(\addr<2> ), .clk(clk), .rst(n1012)
         );
  dff_151 \reg0[3]  ( .q(\addr_1c<3> ), .d(\addr<3> ), .clk(clk), .rst(n1012)
         );
  dff_150 \reg0[4]  ( .q(\addr_1c<4> ), .d(\addr<4> ), .clk(clk), .rst(n1012)
         );
  dff_149 \reg0[5]  ( .q(\addr_1c<5> ), .d(\addr<5> ), .clk(clk), .rst(n1012)
         );
  dff_148 \reg0[6]  ( .q(\addr_1c<6> ), .d(\addr<6> ), .clk(clk), .rst(n1012)
         );
  dff_147 \reg0[7]  ( .q(\addr_1c<7> ), .d(\addr<7> ), .clk(clk), .rst(n1012)
         );
  dff_146 \reg0[8]  ( .q(\addr_1c<8> ), .d(\addr<8> ), .clk(clk), .rst(n1012)
         );
  dff_145 \reg0[9]  ( .q(\addr_1c<9> ), .d(\addr<9> ), .clk(clk), .rst(n1012)
         );
  dff_144 \reg0[10]  ( .q(\addr_1c<10> ), .d(\addr<10> ), .clk(clk), .rst(
        n1012) );
  dff_143 \reg0[11]  ( .q(\addr_1c<11> ), .d(\addr<11> ), .clk(clk), .rst(
        n1012) );
  dff_142 \reg0[12]  ( .q(\addr_1c<12> ), .d(\addr<12> ), .clk(clk), .rst(
        n1012) );
  dff_141 \reg1[0]  ( .q(\data_in_1c<0> ), .d(\data_in<0> ), .clk(clk), .rst(
        n1012) );
  dff_140 \reg1[1]  ( .q(\data_in_1c<1> ), .d(\data_in<1> ), .clk(clk), .rst(
        n1012) );
  dff_139 \reg1[2]  ( .q(\data_in_1c<2> ), .d(\data_in<2> ), .clk(clk), .rst(
        n1012) );
  dff_138 \reg1[3]  ( .q(\data_in_1c<3> ), .d(\data_in<3> ), .clk(clk), .rst(
        n1012) );
  dff_137 \reg1[4]  ( .q(\data_in_1c<4> ), .d(\data_in<4> ), .clk(clk), .rst(
        n1012) );
  dff_136 \reg1[5]  ( .q(\data_in_1c<5> ), .d(\data_in<5> ), .clk(clk), .rst(
        n1012) );
  dff_135 \reg1[6]  ( .q(\data_in_1c<6> ), .d(\data_in<6> ), .clk(clk), .rst(
        n1012) );
  dff_134 \reg1[7]  ( .q(\data_in_1c<7> ), .d(\data_in<7> ), .clk(clk), .rst(
        n1012) );
  dff_133 \reg1[8]  ( .q(\data_in_1c<8> ), .d(\data_in<8> ), .clk(clk), .rst(
        n1012) );
  dff_132 \reg1[9]  ( .q(\data_in_1c<9> ), .d(\data_in<9> ), .clk(clk), .rst(
        n1012) );
  dff_131 \reg1[10]  ( .q(\data_in_1c<10> ), .d(\data_in<10> ), .clk(clk), 
        .rst(n1012) );
  dff_130 \reg1[11]  ( .q(\data_in_1c<11> ), .d(\data_in<11> ), .clk(clk), 
        .rst(n1012) );
  dff_129 \reg1[12]  ( .q(\data_in_1c<12> ), .d(\data_in<12> ), .clk(clk), 
        .rst(n1012) );
  dff_128 \reg1[13]  ( .q(\data_in_1c<13> ), .d(\data_in<13> ), .clk(clk), 
        .rst(n1012) );
  dff_127 \reg1[14]  ( .q(\data_in_1c<14> ), .d(\data_in<14> ), .clk(clk), 
        .rst(n1012) );
  dff_126 \reg1[15]  ( .q(\data_in_1c<15> ), .d(\data_in<15> ), .clk(clk), 
        .rst(n1012) );
  dff_125 \reg2[0]  ( .q(\data_out<0> ), .d(n1022), .clk(clk), .rst(n1012) );
  dff_124 \reg2[1]  ( .q(\data_out<1> ), .d(n1021), .clk(clk), .rst(n1012) );
  dff_123 \reg2[2]  ( .q(\data_out<2> ), .d(n1020), .clk(clk), .rst(n1012) );
  dff_122 \reg2[3]  ( .q(\data_out<3> ), .d(n1019), .clk(clk), .rst(n1012) );
  dff_121 \reg2[4]  ( .q(\data_out<4> ), .d(n1018), .clk(clk), .rst(n1012) );
  dff_120 \reg2[5]  ( .q(\data_out<5> ), .d(n1017), .clk(clk), .rst(n1012) );
  dff_119 \reg2[6]  ( .q(\data_out<6> ), .d(n1016), .clk(clk), .rst(n1012) );
  dff_118 \reg2[7]  ( .q(\data_out<7> ), .d(n1015), .clk(clk), .rst(n1012) );
  dff_117 \reg2[8]  ( .q(\data_out<8> ), .d(\data_out_1c<8> ), .clk(clk), 
        .rst(n1012) );
  dff_116 \reg2[9]  ( .q(\data_out<9> ), .d(\data_out_1c<9> ), .clk(clk), 
        .rst(n1012) );
  dff_115 \reg2[10]  ( .q(\data_out<10> ), .d(\data_out_1c<10> ), .clk(clk), 
        .rst(n1012) );
  dff_114 \reg2[11]  ( .q(\data_out<11> ), .d(\data_out_1c<11> ), .clk(clk), 
        .rst(n1012) );
  dff_113 \reg2[12]  ( .q(\data_out<12> ), .d(\data_out_1c<12> ), .clk(clk), 
        .rst(n1012) );
  dff_112 \reg2[13]  ( .q(\data_out<13> ), .d(\data_out_1c<13> ), .clk(clk), 
        .rst(n1012) );
  dff_111 \reg2[14]  ( .q(\data_out<14> ), .d(\data_out_1c<14> ), .clk(clk), 
        .rst(n1012) );
  dff_110 \reg2[15]  ( .q(\data_out<15> ), .d(\data_out_1c<15> ), .clk(clk), 
        .rst(n1012) );
  dff_109 ff2 ( .q(rd2), .d(rd1), .clk(clk), .rst(n1012) );
  dff_108 ff3 ( .q(wr2), .d(wr1), .clk(clk), .rst(n1012) );
  dff_107 ff4 ( .q(rd3), .d(rd2), .clk(clk), .rst(n1012) );
  dff_106 ff5 ( .q(wr3), .d(wr2), .clk(clk), .rst(n1012) );
  INVX1 U2 ( .A(rd), .Y(n1045) );
  OR2X1 U3 ( .A(\addr_1c<5> ), .B(\addr_1c<12> ), .Y(n1510) );
  AND2X1 U4 ( .A(\addr_1c<4> ), .B(n1524), .Y(n1827) );
  INVX1 U5 ( .A(\addr_1c<3> ), .Y(n1027) );
  INVX1 U6 ( .A(\addr_1c<2> ), .Y(n1026) );
  INVX1 U7 ( .A(wr1), .Y(n1023) );
  INVX1 U8 ( .A(\addr_1c<1> ), .Y(n1025) );
  OR2X1 U23 ( .A(\addr_1c<9> ), .B(\addr_1c<8> ), .Y(n1511) );
  AND2X1 U24 ( .A(\addr_1c<3> ), .B(\addr_1c<0> ), .Y(n1318) );
  AND2X1 U25 ( .A(\addr_1c<3> ), .B(n1024), .Y(n1317) );
  AND2X1 U26 ( .A(n1630), .B(n964), .Y(n1807) );
  AND2X1 U27 ( .A(n1591), .B(n964), .Y(n1766) );
  AND2X1 U28 ( .A(\addr_1c<0> ), .B(n1027), .Y(n1311) );
  AND2X1 U29 ( .A(n1024), .B(n1027), .Y(n1310) );
  INVX1 U35 ( .A(\addr_1c<0> ), .Y(n1024) );
  AND2X1 U36 ( .A(\addr_1c<2> ), .B(n1025), .Y(n1591) );
  AND2X1 U37 ( .A(\addr_1c<2> ), .B(\addr_1c<1> ), .Y(n1630) );
  AND2X1 U38 ( .A(n1317), .B(n1630), .Y(n1796) );
  AND2X1 U39 ( .A(n1591), .B(n1318), .Y(n1776) );
  AND2X1 U40 ( .A(n1591), .B(n1317), .Y(n1756) );
  AND2X1 U41 ( .A(n940), .B(n1318), .Y(n1737) );
  AND2X1 U42 ( .A(n940), .B(n1317), .Y(n1718) );
  AND2X1 U43 ( .A(n1318), .B(n951), .Y(n1699) );
  AND2X1 U44 ( .A(n1317), .B(n951), .Y(n1680) );
  AND2X1 U46 ( .A(n1311), .B(n1630), .Y(n1661) );
  AND2X1 U47 ( .A(n1630), .B(n1310), .Y(n1641) );
  AND2X1 U48 ( .A(n1311), .B(n1591), .Y(n1620) );
  AND2X1 U49 ( .A(n1591), .B(n1310), .Y(n1601) );
  AND2X1 U50 ( .A(n1311), .B(n940), .Y(n1581) );
  AND2X1 U51 ( .A(n940), .B(n1310), .Y(n1562) );
  OR2X1 U52 ( .A(n970), .B(n965), .Y(n968) );
  AND2X1 U53 ( .A(n1311), .B(n951), .Y(n1542) );
  OR2X1 U54 ( .A(n965), .B(n971), .Y(n966) );
  AND2X1 U55 ( .A(n1827), .B(\mem<32><0> ), .Y(n1491) );
  AND2X1 U56 ( .A(n1827), .B(\mem<32><1> ), .Y(n1503) );
  AND2X1 U57 ( .A(n1827), .B(\mem<32><2> ), .Y(n1336) );
  AND2X1 U58 ( .A(n1827), .B(\mem<32><3> ), .Y(n1349) );
  AND2X1 U59 ( .A(n1827), .B(\mem<32><4> ), .Y(n1362) );
  AND2X1 U60 ( .A(n1827), .B(\mem<32><5> ), .Y(n1375) );
  AND2X1 U61 ( .A(n1827), .B(\mem<32><6> ), .Y(n1388) );
  AND2X1 U62 ( .A(n1827), .B(\mem<32><7> ), .Y(n1401) );
  INVX1 U63 ( .A(rd1), .Y(n1014) );
  BUFX2 U64 ( .A(n961), .Y(n1010) );
  BUFX2 U65 ( .A(n961), .Y(n1009) );
  BUFX2 U66 ( .A(n960), .Y(n1007) );
  BUFX2 U67 ( .A(n960), .Y(n1006) );
  BUFX2 U68 ( .A(n959), .Y(n1004) );
  BUFX2 U69 ( .A(n959), .Y(n1003) );
  BUFX2 U70 ( .A(n958), .Y(n1001) );
  BUFX2 U71 ( .A(n958), .Y(n1000) );
  BUFX2 U72 ( .A(n957), .Y(n990) );
  BUFX2 U73 ( .A(n957), .Y(n989) );
  BUFX2 U74 ( .A(n956), .Y(n987) );
  BUFX2 U75 ( .A(n956), .Y(n986) );
  BUFX2 U76 ( .A(n955), .Y(n984) );
  BUFX2 U77 ( .A(n955), .Y(n983) );
  BUFX2 U78 ( .A(n954), .Y(n981) );
  BUFX2 U79 ( .A(n954), .Y(n980) );
  INVX1 U80 ( .A(\data_in_1c<0> ), .Y(n1028) );
  INVX1 U81 ( .A(\data_in_1c<1> ), .Y(n1029) );
  INVX1 U82 ( .A(\data_in_1c<2> ), .Y(n1030) );
  INVX1 U83 ( .A(\data_in_1c<3> ), .Y(n1031) );
  INVX1 U84 ( .A(\data_in_1c<4> ), .Y(n1032) );
  INVX1 U85 ( .A(\data_in_1c<5> ), .Y(n1033) );
  INVX1 U86 ( .A(\data_in_1c<6> ), .Y(n1034) );
  INVX1 U87 ( .A(\data_in_1c<7> ), .Y(n1035) );
  INVX1 U88 ( .A(\data_in_1c<8> ), .Y(n1036) );
  INVX1 U89 ( .A(\data_in_1c<9> ), .Y(n1037) );
  INVX1 U90 ( .A(\data_in_1c<10> ), .Y(n1038) );
  INVX1 U91 ( .A(\data_in_1c<11> ), .Y(n1039) );
  INVX1 U92 ( .A(\data_in_1c<12> ), .Y(n1040) );
  INVX1 U93 ( .A(\data_in_1c<13> ), .Y(n1041) );
  INVX1 U129 ( .A(\data_in_1c<14> ), .Y(n1042) );
  INVX1 U589 ( .A(\data_in_1c<15> ), .Y(n1043) );
  INVX1 U640 ( .A(wr), .Y(n1044) );
  INVX1 U659 ( .A(n1324), .Y(n1022) );
  INVX1 U660 ( .A(n1415), .Y(n1021) );
  INVX1 U664 ( .A(n1426), .Y(n1020) );
  INVX1 U666 ( .A(n1437), .Y(n1019) );
  INVX1 U672 ( .A(n1448), .Y(n1018) );
  INVX1 U675 ( .A(n1459), .Y(n1017) );
  INVX1 U679 ( .A(n1470), .Y(n1016) );
  INVX1 U682 ( .A(n1481), .Y(n1015) );
  INVX1 U694 ( .A(rst), .Y(n1013) );
  INVX2 U697 ( .A(n1013), .Y(n1012) );
  AND2X1 U701 ( .A(wr1), .B(n1013), .Y(n1828) );
  AND2X1 U706 ( .A(n387), .B(n372), .Y(n1) );
  INVX1 U712 ( .A(n1), .Y(n2) );
  AND2X1 U717 ( .A(n402), .B(n381), .Y(n3) );
  INVX1 U723 ( .A(n3), .Y(n4) );
  AND2X1 U728 ( .A(n1817), .B(n189), .Y(n5) );
  INVX1 U734 ( .A(n5), .Y(n6) );
  AND2X1 U739 ( .A(n973), .B(n289), .Y(n7) );
  INVX1 U745 ( .A(n7), .Y(n8) );
  OR2X1 U750 ( .A(n486), .B(n10), .Y(n9) );
  OR2X1 U756 ( .A(n473), .B(n474), .Y(n10) );
  OR2X1 U761 ( .A(n508), .B(n12), .Y(n11) );
  OR2X1 U767 ( .A(n487), .B(n507), .Y(n12) );
  OR2X1 U772 ( .A(n537), .B(n14), .Y(n13) );
  OR2X1 U786 ( .A(n522), .B(n523), .Y(n14) );
  OR2X1 U789 ( .A(n553), .B(n16), .Y(n15) );
  OR2X1 U801 ( .A(n538), .B(n552), .Y(n16) );
  OR2X1 U804 ( .A(n582), .B(n18), .Y(n17) );
  OR2X1 U816 ( .A(n567), .B(n568), .Y(n18) );
  OR2X1 U819 ( .A(n592), .B(n20), .Y(n19) );
  OR2X1 U831 ( .A(n583), .B(n591), .Y(n20) );
  OR2X1 U834 ( .A(n873), .B(n22), .Y(n21) );
  OR2X1 U846 ( .A(n871), .B(n872), .Y(n22) );
  OR2X1 U849 ( .A(n876), .B(n24), .Y(n23) );
  OR2X1 U861 ( .A(n874), .B(n875), .Y(n24) );
  OR2X1 U864 ( .A(n895), .B(n26), .Y(n25) );
  OR2X1 U870 ( .A(n893), .B(n894), .Y(n26) );
  OR2X1 U875 ( .A(n898), .B(n28), .Y(n27) );
  OR2X1 U882 ( .A(n896), .B(n897), .Y(n28) );
  OR2X1 U883 ( .A(n901), .B(n30), .Y(n29) );
  OR2X1 U884 ( .A(n899), .B(n900), .Y(n30) );
  OR2X1 U885 ( .A(n904), .B(n32), .Y(n31) );
  OR2X1 U886 ( .A(n902), .B(n903), .Y(n32) );
  OR2X1 U887 ( .A(n907), .B(n34), .Y(n33) );
  OR2X1 U888 ( .A(n905), .B(n906), .Y(n34) );
  OR2X1 U889 ( .A(n910), .B(n36), .Y(n35) );
  OR2X1 U890 ( .A(n908), .B(n909), .Y(n36) );
  OR2X1 U891 ( .A(n913), .B(n38), .Y(n37) );
  OR2X1 U892 ( .A(n911), .B(n912), .Y(n38) );
  OR2X1 U893 ( .A(n916), .B(n150), .Y(n50) );
  OR2X1 U894 ( .A(n914), .B(n915), .Y(n150) );
  AND2X1 U895 ( .A(n973), .B(n1828), .Y(n189) );
  AND2X1 U896 ( .A(n1828), .B(n1524), .Y(n289) );
  AND2X1 U897 ( .A(n940), .B(n942), .Y(n348) );
  INVX1 U898 ( .A(n348), .Y(n372) );
  AND2X1 U899 ( .A(n951), .B(n953), .Y(n379) );
  INVX1 U900 ( .A(n379), .Y(n381) );
  AND2X1 U901 ( .A(n940), .B(n941), .Y(n386) );
  INVX1 U902 ( .A(n386), .Y(n387) );
  AND2X1 U903 ( .A(n951), .B(n952), .Y(n401) );
  INVX1 U904 ( .A(n401), .Y(n402) );
  BUFX2 U905 ( .A(n1339), .Y(n408) );
  BUFX2 U906 ( .A(n1352), .Y(n409) );
  BUFX2 U907 ( .A(n1365), .Y(n421) );
  BUFX2 U908 ( .A(n1378), .Y(n422) );
  BUFX2 U909 ( .A(n1391), .Y(n434) );
  BUFX2 U910 ( .A(n1404), .Y(n435) );
  BUFX2 U911 ( .A(n1494), .Y(n447) );
  BUFX2 U912 ( .A(n1505), .Y(n448) );
  AND2X2 U913 ( .A(rd), .B(n1508), .Y(n460) );
  INVX1 U914 ( .A(n460), .Y(n461) );
  INVX1 U915 ( .A(n1314), .Y(n473) );
  INVX1 U916 ( .A(n1315), .Y(n474) );
  INVX1 U917 ( .A(n1316), .Y(n486) );
  INVX1 U918 ( .A(n1407), .Y(n487) );
  INVX1 U919 ( .A(n1408), .Y(n507) );
  INVX1 U920 ( .A(n1409), .Y(n508) );
  INVX1 U921 ( .A(n1418), .Y(n522) );
  INVX1 U922 ( .A(n1419), .Y(n523) );
  INVX1 U923 ( .A(n1420), .Y(n537) );
  INVX1 U924 ( .A(n1429), .Y(n538) );
  INVX1 U925 ( .A(n1430), .Y(n552) );
  INVX1 U926 ( .A(n1431), .Y(n553) );
  INVX1 U927 ( .A(n1440), .Y(n567) );
  INVX1 U928 ( .A(n1441), .Y(n568) );
  INVX1 U929 ( .A(n1442), .Y(n582) );
  INVX1 U930 ( .A(n1451), .Y(n583) );
  INVX1 U931 ( .A(n1452), .Y(n591) );
  INVX1 U932 ( .A(n1453), .Y(n592) );
  INVX1 U933 ( .A(n1462), .Y(n871) );
  INVX1 U934 ( .A(n1463), .Y(n872) );
  INVX1 U935 ( .A(n1464), .Y(n873) );
  INVX1 U936 ( .A(n1473), .Y(n874) );
  INVX1 U937 ( .A(n1474), .Y(n875) );
  INVX1 U938 ( .A(n1475), .Y(n876) );
  AND2X2 U939 ( .A(n1328), .B(n1327), .Y(n877) );
  INVX1 U940 ( .A(n877), .Y(n878) );
  AND2X2 U941 ( .A(n1341), .B(n1340), .Y(n879) );
  INVX1 U942 ( .A(n879), .Y(n880) );
  AND2X2 U943 ( .A(n1354), .B(n1353), .Y(n881) );
  INVX1 U944 ( .A(n881), .Y(n882) );
  AND2X2 U945 ( .A(n1367), .B(n1366), .Y(n883) );
  INVX1 U946 ( .A(n883), .Y(n884) );
  AND2X2 U947 ( .A(n1380), .B(n1379), .Y(n885) );
  INVX1 U948 ( .A(n885), .Y(n886) );
  AND2X2 U949 ( .A(n1393), .B(n1392), .Y(n887) );
  INVX1 U950 ( .A(n887), .Y(n888) );
  AND2X2 U951 ( .A(n1483), .B(n1482), .Y(n889) );
  INVX1 U952 ( .A(n889), .Y(n890) );
  AND2X2 U953 ( .A(n1496), .B(n1495), .Y(n891) );
  INVX1 U954 ( .A(n891), .Y(n892) );
  INVX1 U955 ( .A(n1321), .Y(n893) );
  INVX1 U956 ( .A(n1322), .Y(n894) );
  INVX1 U957 ( .A(n1323), .Y(n895) );
  INVX1 U958 ( .A(n1412), .Y(n896) );
  INVX1 U959 ( .A(n1413), .Y(n897) );
  INVX1 U960 ( .A(n1414), .Y(n898) );
  INVX1 U961 ( .A(n1423), .Y(n899) );
  INVX1 U962 ( .A(n1424), .Y(n900) );
  INVX1 U963 ( .A(n1425), .Y(n901) );
  INVX1 U964 ( .A(n1434), .Y(n902) );
  INVX1 U965 ( .A(n1435), .Y(n903) );
  INVX1 U966 ( .A(n1436), .Y(n904) );
  INVX1 U967 ( .A(n1445), .Y(n905) );
  INVX1 U968 ( .A(n1446), .Y(n906) );
  INVX1 U969 ( .A(n1447), .Y(n907) );
  INVX1 U970 ( .A(n1456), .Y(n908) );
  INVX1 U971 ( .A(n1457), .Y(n909) );
  INVX1 U972 ( .A(n1458), .Y(n910) );
  INVX1 U973 ( .A(n1467), .Y(n911) );
  INVX1 U974 ( .A(n1468), .Y(n912) );
  INVX1 U975 ( .A(n1469), .Y(n913) );
  INVX1 U976 ( .A(n1478), .Y(n914) );
  INVX1 U977 ( .A(n1479), .Y(n915) );
  INVX1 U978 ( .A(n1480), .Y(n916) );
  AND2X2 U979 ( .A(n1330), .B(n1329), .Y(n917) );
  INVX1 U980 ( .A(n917), .Y(n918) );
  AND2X2 U981 ( .A(n1343), .B(n1342), .Y(n919) );
  INVX1 U982 ( .A(n919), .Y(n920) );
  AND2X2 U983 ( .A(n1356), .B(n1355), .Y(n921) );
  INVX1 U984 ( .A(n921), .Y(n922) );
  AND2X2 U985 ( .A(n1369), .B(n1368), .Y(n923) );
  INVX1 U986 ( .A(n923), .Y(n924) );
  AND2X2 U987 ( .A(n1382), .B(n1381), .Y(n925) );
  INVX1 U988 ( .A(n925), .Y(n926) );
  AND2X2 U989 ( .A(n1395), .B(n1394), .Y(n927) );
  INVX1 U990 ( .A(n927), .Y(n928) );
  AND2X2 U991 ( .A(n1485), .B(n1484), .Y(n929) );
  INVX1 U992 ( .A(n929), .Y(n930) );
  AND2X2 U993 ( .A(n1498), .B(n1497), .Y(n931) );
  INVX1 U994 ( .A(n931), .Y(n932) );
  BUFX2 U995 ( .A(n1337), .Y(n933) );
  BUFX2 U996 ( .A(n1350), .Y(n934) );
  BUFX2 U997 ( .A(n1363), .Y(n935) );
  BUFX2 U998 ( .A(n1376), .Y(n936) );
  BUFX2 U999 ( .A(n1389), .Y(n937) );
  BUFX2 U1000 ( .A(n1402), .Y(n938) );
  BUFX2 U1001 ( .A(n1492), .Y(n939) );
  INVX1 U1002 ( .A(n970), .Y(n940) );
  INVX1 U1003 ( .A(n1499), .Y(n941) );
  INVX1 U1004 ( .A(n1500), .Y(n942) );
  BUFX2 U1005 ( .A(n1552), .Y(n970) );
  BUFX2 U1006 ( .A(n1838), .Y(err) );
  BUFX2 U1007 ( .A(n1335), .Y(n944) );
  BUFX2 U1008 ( .A(n1348), .Y(n945) );
  BUFX2 U1009 ( .A(n1361), .Y(n946) );
  BUFX2 U1010 ( .A(n1374), .Y(n947) );
  BUFX2 U1011 ( .A(n1387), .Y(n948) );
  BUFX2 U1012 ( .A(n1400), .Y(n949) );
  BUFX2 U1013 ( .A(n1490), .Y(n950) );
  INVX1 U1014 ( .A(n971), .Y(n951) );
  INVX1 U1015 ( .A(n1501), .Y(n952) );
  INVX1 U1016 ( .A(n1502), .Y(n953) );
  BUFX2 U1017 ( .A(n1514), .Y(n971) );
  BUFX2 U1018 ( .A(n1523), .Y(n972) );
  BUFX2 U1019 ( .A(n1541), .Y(n974) );
  BUFX2 U1020 ( .A(n1551), .Y(n975) );
  BUFX2 U1021 ( .A(n1561), .Y(n976) );
  BUFX2 U1022 ( .A(n1571), .Y(n977) );
  BUFX2 U1023 ( .A(n1580), .Y(n978) );
  BUFX2 U1024 ( .A(n1590), .Y(n979) );
  BUFX2 U1025 ( .A(n1610), .Y(n982) );
  BUFX2 U1026 ( .A(n1629), .Y(n985) );
  BUFX2 U1027 ( .A(n1650), .Y(n988) );
  BUFX2 U1028 ( .A(n1670), .Y(n991) );
  BUFX2 U1029 ( .A(n1679), .Y(n992) );
  BUFX2 U1030 ( .A(n1689), .Y(n993) );
  BUFX2 U1031 ( .A(n1698), .Y(n994) );
  BUFX2 U1032 ( .A(n1708), .Y(n995) );
  BUFX2 U1033 ( .A(n1717), .Y(n996) );
  BUFX2 U1034 ( .A(n1727), .Y(n997) );
  BUFX2 U1035 ( .A(n1736), .Y(n998) );
  BUFX2 U1036 ( .A(n1746), .Y(n999) );
  BUFX2 U1037 ( .A(n1765), .Y(n1002) );
  BUFX2 U1038 ( .A(n1785), .Y(n1005) );
  BUFX2 U1039 ( .A(n1805), .Y(n1008) );
  BUFX2 U1040 ( .A(n1818), .Y(n973) );
  AND2X1 U1041 ( .A(n1630), .B(n1318), .Y(n1817) );
  BUFX2 U1042 ( .A(n1837), .Y(n1011) );
  BUFX2 U1043 ( .A(n1600), .Y(n954) );
  BUFX2 U1044 ( .A(n1619), .Y(n955) );
  BUFX2 U1045 ( .A(n1640), .Y(n956) );
  BUFX2 U1046 ( .A(n1660), .Y(n957) );
  BUFX2 U1047 ( .A(n1755), .Y(n958) );
  BUFX2 U1048 ( .A(n1775), .Y(n959) );
  BUFX2 U1049 ( .A(n1795), .Y(n960) );
  BUFX2 U1050 ( .A(n1816), .Y(n961) );
  AND2X1 U1051 ( .A(enable), .B(n1013), .Y(n962) );
  INVX1 U1052 ( .A(n962), .Y(n963) );
  AND2X1 U1053 ( .A(n1513), .B(n1512), .Y(n964) );
  INVX1 U1054 ( .A(n964), .Y(n965) );
  INVX1 U1055 ( .A(n966), .Y(n967) );
  INVX1 U1056 ( .A(n968), .Y(n969) );
  AND2X1 U1057 ( .A(n951), .B(n1310), .Y(n1524) );
endmodule


module final_memory_1 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), err, .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<12> , \addr<11> , \addr<10> , \addr<9> , 
        \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , 
        \addr<2> , \addr<1> , \addr<0> }), wr, rd, enable, create_dump, 
    .bank_id({\bank_id<1> , \bank_id<0> }), clk, rst );
  input \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , \addr<12> , \addr<11> ,
         \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> , \addr<5> ,
         \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> , wr, rd, enable,
         create_dump, \bank_id<1> , \bank_id<0> , clk, rst;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , err;
  wire   n1838, rd0, wr0, rd1, wr1, \addr_1c<12> , \addr_1c<11> ,
         \addr_1c<10> , \addr_1c<9> , \addr_1c<8> , \addr_1c<7> , \addr_1c<6> ,
         \addr_1c<5> , \addr_1c<4> , \addr_1c<3> , \addr_1c<2> , \addr_1c<1> ,
         \addr_1c<0> , \data_in_1c<15> , \data_in_1c<14> , \data_in_1c<13> ,
         \data_in_1c<12> , \data_in_1c<11> , \data_in_1c<10> , \data_in_1c<9> ,
         \data_in_1c<8> , \data_in_1c<7> , \data_in_1c<6> , \data_in_1c<5> ,
         \data_in_1c<4> , \data_in_1c<3> , \data_in_1c<2> , \data_in_1c<1> ,
         \data_in_1c<0> , \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> ,
         \mem<0><3> , \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><7> ,
         \mem<1><6> , \mem<1><5> , \mem<1><4> , \mem<1><3> , \mem<1><2> ,
         \mem<1><1> , \mem<1><0> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><7> , \mem<3><6> , \mem<3><5> , \mem<3><4> , \mem<3><3> ,
         \mem<3><2> , \mem<3><1> , \mem<3><0> , \mem<4><7> , \mem<4><6> ,
         \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> , \mem<4><1> ,
         \mem<4><0> , \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> ,
         \mem<5><3> , \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><7> ,
         \mem<6><6> , \mem<6><5> , \mem<6><4> , \mem<6><3> , \mem<6><2> ,
         \mem<6><1> , \mem<6><0> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><7> , \mem<8><6> , \mem<8><5> , \mem<8><4> , \mem<8><3> ,
         \mem<8><2> , \mem<8><1> , \mem<8><0> , \mem<9><7> , \mem<9><6> ,
         \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> , \mem<9><1> ,
         \mem<9><0> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><7> ,
         \mem<11><6> , \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> ,
         \mem<11><1> , \mem<11><0> , \mem<12><7> , \mem<12><6> , \mem<12><5> ,
         \mem<12><4> , \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> ,
         \mem<13><7> , \mem<13><6> , \mem<13><5> , \mem<13><4> , \mem<13><3> ,
         \mem<13><2> , \mem<13><1> , \mem<13><0> , \mem<14><7> , \mem<14><6> ,
         \mem<14><5> , \mem<14><4> , \mem<14><3> , \mem<14><2> , \mem<14><1> ,
         \mem<14><0> , \mem<15><7> , \mem<15><6> , \mem<15><5> , \mem<15><4> ,
         \mem<15><3> , \mem<15><2> , \mem<15><1> , \mem<15><0> , \mem<16><7> ,
         \mem<16><6> , \mem<16><5> , \mem<16><4> , \mem<16><3> , \mem<16><2> ,
         \mem<16><1> , \mem<16><0> , \mem<17><7> , \mem<17><6> , \mem<17><5> ,
         \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> , \mem<17><0> ,
         \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> , \mem<18><3> ,
         \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><7> ,
         \mem<21><6> , \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> ,
         \mem<21><1> , \mem<21><0> , \mem<22><7> , \mem<22><6> , \mem<22><5> ,
         \mem<22><4> , \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> ,
         \mem<23><7> , \mem<23><6> , \mem<23><5> , \mem<23><4> , \mem<23><3> ,
         \mem<23><2> , \mem<23><1> , \mem<23><0> , \mem<24><7> , \mem<24><6> ,
         \mem<24><5> , \mem<24><4> , \mem<24><3> , \mem<24><2> , \mem<24><1> ,
         \mem<24><0> , \mem<25><7> , \mem<25><6> , \mem<25><5> , \mem<25><4> ,
         \mem<25><3> , \mem<25><2> , \mem<25><1> , \mem<25><0> , \mem<26><7> ,
         \mem<26><6> , \mem<26><5> , \mem<26><4> , \mem<26><3> , \mem<26><2> ,
         \mem<26><1> , \mem<26><0> , \mem<27><7> , \mem<27><6> , \mem<27><5> ,
         \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> , \mem<27><0> ,
         \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> , \mem<28><3> ,
         \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><7> ,
         \mem<31><6> , \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> ,
         \mem<31><1> , \mem<31><0> , \mem<32><7> , \mem<32><6> , \mem<32><5> ,
         \mem<32><4> , \mem<32><3> , \mem<32><2> , \mem<32><1> , \mem<32><0> ,
         \data_out_1c<15> , \data_out_1c<14> , \data_out_1c<13> ,
         \data_out_1c<12> , \data_out_1c<11> , \data_out_1c<10> ,
         \data_out_1c<9> , \data_out_1c<8> , rd2, wr2, rd3, wr3, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n50, n150, n189, n289, n348, n372, n379,
         n381, n386, n387, n401, n402, n408, n409, n421, n422, n434, n435,
         n447, n448, n460, n461, n473, n474, n486, n487, n507, n508, n522,
         n523, n537, n538, n552, n553, n567, n568, n582, n583, n591, n592,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837;

  DFFPOSX1 \mem_reg<0><7>  ( .D(n1046), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1047), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1048), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1049), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1050), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1051), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1052), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1053), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1054), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1055), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1056), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1057), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1058), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1059), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1060), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1061), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1062), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1063), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1064), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1065), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1066), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1067), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1068), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1069), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1070), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1071), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1072), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1073), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1074), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1075), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1076), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1077), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1078), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1079), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1080), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1081), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1082), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1083), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1084), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1085), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1086), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1087), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1088), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1089), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1090), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1091), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1092), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1093), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1094), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1095), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1096), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1097), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1098), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1099), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1100), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1101), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1102), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1103), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1104), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1105), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1106), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1107), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1108), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1109), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1110), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1111), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1112), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1113), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1114), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1115), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1116), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1117), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n1118), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n1119), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n1120), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n1121), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n1122), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n1123), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n1124), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n1125), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n1126), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n1127), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n1128), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n1129), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n1130), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n1131), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n1132), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n1133), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n1134), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n1135), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n1136), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n1137), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n1138), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n1139), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n1140), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n1141), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n1142), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n1143), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n1144), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n1145), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n1146), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n1147), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n1148), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n1149), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n1150), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n1151), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n1152), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n1153), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n1154), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n1155), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n1156), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n1157), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n1158), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n1159), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n1160), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n1161), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n1162), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n1163), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n1164), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n1165), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n1166), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n1167), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n1168), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n1169), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n1170), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n1171), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n1172), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n1173), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n1174), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n1175), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n1176), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n1177), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n1178), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n1179), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n1180), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n1181), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n1182), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n1183), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n1184), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n1185), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n1186), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n1187), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n1188), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n1189), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n1190), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n1191), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n1192), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n1193), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n1194), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n1195), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n1196), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n1197), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n1198), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n1199), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n1200), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n1201), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n1202), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n1203), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n1204), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n1205), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n1206), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n1207), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n1208), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n1209), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n1210), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n1211), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n1212), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n1213), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n1214), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n1215), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n1216), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n1217), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n1218), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n1219), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n1220), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n1221), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n1222), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n1223), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n1224), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n1225), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n1226), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n1227), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n1228), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n1229), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n1230), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n1231), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n1232), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n1233), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n1234), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n1235), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n1236), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n1237), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n1238), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n1239), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n1240), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n1241), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n1242), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n1243), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n1244), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n1245), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n1246), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n1247), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n1248), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n1249), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n1250), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n1251), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n1252), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n1253), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n1254), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n1255), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n1256), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n1257), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n1258), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n1259), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n1260), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n1261), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n1262), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n1263), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n1264), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n1265), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n1266), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n1267), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n1268), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n1269), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n1270), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n1271), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n1272), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n1273), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n1274), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n1275), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n1276), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n1277), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n1278), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n1279), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n1280), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n1281), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n1282), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n1283), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n1284), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n1285), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n1286), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n1287), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n1288), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n1289), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n1290), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n1291), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n1292), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n1293), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n1294), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n1295), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n1296), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n1297), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n1298), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n1299), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n1300), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n1301), .CLK(clk), .Q(\mem<31><0> ) );
  DFFPOSX1 \mem_reg<32><7>  ( .D(n1302), .CLK(clk), .Q(\mem<32><7> ) );
  DFFPOSX1 \mem_reg<32><6>  ( .D(n1303), .CLK(clk), .Q(\mem<32><6> ) );
  DFFPOSX1 \mem_reg<32><5>  ( .D(n1304), .CLK(clk), .Q(\mem<32><5> ) );
  DFFPOSX1 \mem_reg<32><4>  ( .D(n1305), .CLK(clk), .Q(\mem<32><4> ) );
  DFFPOSX1 \mem_reg<32><3>  ( .D(n1306), .CLK(clk), .Q(\mem<32><3> ) );
  DFFPOSX1 \mem_reg<32><2>  ( .D(n1307), .CLK(clk), .Q(\mem<32><2> ) );
  DFFPOSX1 \mem_reg<32><1>  ( .D(n1308), .CLK(clk), .Q(\mem<32><1> ) );
  DFFPOSX1 \mem_reg<32><0>  ( .D(n1309), .CLK(clk), .Q(\mem<32><0> ) );
  AND2X2 U9 ( .A(n1477), .B(n1476), .Y(n1478) );
  AND2X2 U10 ( .A(n1472), .B(n1471), .Y(n1473) );
  AND2X2 U11 ( .A(n1466), .B(n1465), .Y(n1467) );
  AND2X2 U12 ( .A(n1461), .B(n1460), .Y(n1462) );
  AND2X2 U13 ( .A(n1455), .B(n1454), .Y(n1456) );
  AND2X2 U14 ( .A(n1450), .B(n1449), .Y(n1451) );
  AND2X2 U15 ( .A(n1444), .B(n1443), .Y(n1445) );
  AND2X2 U16 ( .A(n1439), .B(n1438), .Y(n1440) );
  AND2X2 U17 ( .A(n1433), .B(n1432), .Y(n1434) );
  AND2X2 U18 ( .A(n1428), .B(n1427), .Y(n1429) );
  AND2X2 U19 ( .A(n1422), .B(n1421), .Y(n1423) );
  AND2X2 U20 ( .A(n1417), .B(n1416), .Y(n1418) );
  AND2X2 U21 ( .A(n1411), .B(n1410), .Y(n1412) );
  AND2X2 U22 ( .A(n1406), .B(n1405), .Y(n1407) );
  AND2X2 U30 ( .A(n1326), .B(n1024), .Y(n1631) );
  AND2X2 U31 ( .A(n1325), .B(n1024), .Y(n1786) );
  AND2X2 U32 ( .A(n1326), .B(\addr_1c<0> ), .Y(n1651) );
  AND2X2 U33 ( .A(n1325), .B(\addr_1c<0> ), .Y(n1806) );
  AND2X2 U34 ( .A(n1320), .B(n1319), .Y(n1321) );
  AND2X2 U45 ( .A(n1313), .B(n1312), .Y(n1314) );
  NOR3X1 U94 ( .A(n1044), .B(rd), .C(n963), .Y(wr0) );
  NOR3X1 U95 ( .A(n1045), .B(wr), .C(n963), .Y(rd0) );
  OAI21X1 U96 ( .A(n1011), .B(n1036), .C(n1836), .Y(n1309) );
  NAND2X1 U97 ( .A(\mem<32><0> ), .B(n1011), .Y(n1836) );
  OAI21X1 U98 ( .A(n1011), .B(n1037), .C(n1835), .Y(n1308) );
  NAND2X1 U99 ( .A(\mem<32><1> ), .B(n1011), .Y(n1835) );
  OAI21X1 U100 ( .A(n1011), .B(n1038), .C(n1834), .Y(n1307) );
  NAND2X1 U101 ( .A(\mem<32><2> ), .B(n1011), .Y(n1834) );
  OAI21X1 U102 ( .A(n1011), .B(n1039), .C(n1833), .Y(n1306) );
  NAND2X1 U103 ( .A(\mem<32><3> ), .B(n1011), .Y(n1833) );
  OAI21X1 U104 ( .A(n1011), .B(n1040), .C(n1832), .Y(n1305) );
  NAND2X1 U105 ( .A(\mem<32><4> ), .B(n1011), .Y(n1832) );
  OAI21X1 U106 ( .A(n1011), .B(n1041), .C(n1831), .Y(n1304) );
  NAND2X1 U107 ( .A(\mem<32><5> ), .B(n1011), .Y(n1831) );
  OAI21X1 U108 ( .A(n1011), .B(n1042), .C(n1830), .Y(n1303) );
  NAND2X1 U109 ( .A(\mem<32><6> ), .B(n1011), .Y(n1830) );
  OAI21X1 U110 ( .A(n1011), .B(n1043), .C(n1829), .Y(n1302) );
  NAND2X1 U111 ( .A(\mem<32><7> ), .B(n1011), .Y(n1829) );
  NAND3X1 U112 ( .A(n1828), .B(n1827), .C(n964), .Y(n1837) );
  OAI21X1 U113 ( .A(n6), .B(n1028), .C(n1826), .Y(n1301) );
  NAND2X1 U114 ( .A(\mem<31><0> ), .B(n6), .Y(n1826) );
  OAI21X1 U115 ( .A(n6), .B(n1029), .C(n1825), .Y(n1300) );
  NAND2X1 U116 ( .A(\mem<31><1> ), .B(n6), .Y(n1825) );
  OAI21X1 U117 ( .A(n6), .B(n1030), .C(n1824), .Y(n1299) );
  NAND2X1 U118 ( .A(\mem<31><2> ), .B(n6), .Y(n1824) );
  OAI21X1 U119 ( .A(n6), .B(n1031), .C(n1823), .Y(n1298) );
  NAND2X1 U120 ( .A(\mem<31><3> ), .B(n6), .Y(n1823) );
  OAI21X1 U121 ( .A(n6), .B(n1032), .C(n1822), .Y(n1297) );
  NAND2X1 U122 ( .A(\mem<31><4> ), .B(n6), .Y(n1822) );
  OAI21X1 U123 ( .A(n6), .B(n1033), .C(n1821), .Y(n1296) );
  NAND2X1 U124 ( .A(\mem<31><5> ), .B(n6), .Y(n1821) );
  OAI21X1 U125 ( .A(n6), .B(n1034), .C(n1820), .Y(n1295) );
  NAND2X1 U126 ( .A(\mem<31><6> ), .B(n6), .Y(n1820) );
  OAI21X1 U127 ( .A(n6), .B(n1035), .C(n1819), .Y(n1294) );
  NAND2X1 U128 ( .A(\mem<31><7> ), .B(n6), .Y(n1819) );
  OAI21X1 U130 ( .A(n1036), .B(n1010), .C(n1815), .Y(n1293) );
  NAND2X1 U131 ( .A(\mem<30><0> ), .B(n1010), .Y(n1815) );
  OAI21X1 U132 ( .A(n1037), .B(n1009), .C(n1814), .Y(n1292) );
  NAND2X1 U133 ( .A(\mem<30><1> ), .B(n1010), .Y(n1814) );
  OAI21X1 U134 ( .A(n1038), .B(n1009), .C(n1813), .Y(n1291) );
  NAND2X1 U135 ( .A(\mem<30><2> ), .B(n1010), .Y(n1813) );
  OAI21X1 U136 ( .A(n1039), .B(n1009), .C(n1812), .Y(n1290) );
  NAND2X1 U137 ( .A(\mem<30><3> ), .B(n1010), .Y(n1812) );
  OAI21X1 U138 ( .A(n1040), .B(n1009), .C(n1811), .Y(n1289) );
  NAND2X1 U139 ( .A(\mem<30><4> ), .B(n1010), .Y(n1811) );
  OAI21X1 U140 ( .A(n1041), .B(n1009), .C(n1810), .Y(n1288) );
  NAND2X1 U141 ( .A(\mem<30><5> ), .B(n1010), .Y(n1810) );
  OAI21X1 U142 ( .A(n1042), .B(n1009), .C(n1809), .Y(n1287) );
  NAND2X1 U143 ( .A(\mem<30><6> ), .B(n1010), .Y(n1809) );
  OAI21X1 U144 ( .A(n1043), .B(n1009), .C(n1808), .Y(n1286) );
  NAND2X1 U145 ( .A(\mem<30><7> ), .B(n1010), .Y(n1808) );
  NAND3X1 U146 ( .A(n1807), .B(n1828), .C(n1806), .Y(n1816) );
  OAI21X1 U147 ( .A(n1028), .B(n1008), .C(n1804), .Y(n1285) );
  NAND2X1 U148 ( .A(\mem<29><0> ), .B(n1008), .Y(n1804) );
  OAI21X1 U149 ( .A(n1029), .B(n1008), .C(n1803), .Y(n1284) );
  NAND2X1 U150 ( .A(\mem<29><1> ), .B(n1008), .Y(n1803) );
  OAI21X1 U151 ( .A(n1030), .B(n1008), .C(n1802), .Y(n1283) );
  NAND2X1 U152 ( .A(\mem<29><2> ), .B(n1008), .Y(n1802) );
  OAI21X1 U153 ( .A(n1031), .B(n1008), .C(n1801), .Y(n1282) );
  NAND2X1 U154 ( .A(\mem<29><3> ), .B(n1008), .Y(n1801) );
  OAI21X1 U155 ( .A(n1032), .B(n1008), .C(n1800), .Y(n1281) );
  NAND2X1 U156 ( .A(\mem<29><4> ), .B(n1008), .Y(n1800) );
  OAI21X1 U157 ( .A(n1033), .B(n1008), .C(n1799), .Y(n1280) );
  NAND2X1 U158 ( .A(\mem<29><5> ), .B(n1008), .Y(n1799) );
  OAI21X1 U159 ( .A(n1034), .B(n1008), .C(n1798), .Y(n1279) );
  NAND2X1 U160 ( .A(\mem<29><6> ), .B(n1008), .Y(n1798) );
  OAI21X1 U161 ( .A(n1035), .B(n1008), .C(n1797), .Y(n1278) );
  NAND2X1 U162 ( .A(\mem<29><7> ), .B(n1008), .Y(n1797) );
  NAND3X1 U163 ( .A(n973), .B(n1828), .C(n1796), .Y(n1805) );
  OAI21X1 U164 ( .A(n1036), .B(n1007), .C(n1794), .Y(n1277) );
  NAND2X1 U165 ( .A(\mem<28><0> ), .B(n1007), .Y(n1794) );
  OAI21X1 U166 ( .A(n1037), .B(n1006), .C(n1793), .Y(n1276) );
  NAND2X1 U167 ( .A(\mem<28><1> ), .B(n1007), .Y(n1793) );
  OAI21X1 U168 ( .A(n1038), .B(n1006), .C(n1792), .Y(n1275) );
  NAND2X1 U169 ( .A(\mem<28><2> ), .B(n1007), .Y(n1792) );
  OAI21X1 U170 ( .A(n1039), .B(n1006), .C(n1791), .Y(n1274) );
  NAND2X1 U171 ( .A(\mem<28><3> ), .B(n1007), .Y(n1791) );
  OAI21X1 U172 ( .A(n1040), .B(n1006), .C(n1790), .Y(n1273) );
  NAND2X1 U173 ( .A(\mem<28><4> ), .B(n1007), .Y(n1790) );
  OAI21X1 U174 ( .A(n1041), .B(n1006), .C(n1789), .Y(n1272) );
  NAND2X1 U175 ( .A(\mem<28><5> ), .B(n1007), .Y(n1789) );
  OAI21X1 U176 ( .A(n1042), .B(n1006), .C(n1788), .Y(n1271) );
  NAND2X1 U177 ( .A(\mem<28><6> ), .B(n1007), .Y(n1788) );
  OAI21X1 U178 ( .A(n1043), .B(n1006), .C(n1787), .Y(n1270) );
  NAND2X1 U179 ( .A(\mem<28><7> ), .B(n1007), .Y(n1787) );
  NAND3X1 U180 ( .A(n1807), .B(n1828), .C(n1786), .Y(n1795) );
  OAI21X1 U181 ( .A(n1028), .B(n1005), .C(n1784), .Y(n1269) );
  NAND2X1 U182 ( .A(\mem<27><0> ), .B(n1005), .Y(n1784) );
  OAI21X1 U183 ( .A(n1029), .B(n1005), .C(n1783), .Y(n1268) );
  NAND2X1 U184 ( .A(\mem<27><1> ), .B(n1005), .Y(n1783) );
  OAI21X1 U185 ( .A(n1030), .B(n1005), .C(n1782), .Y(n1267) );
  NAND2X1 U186 ( .A(\mem<27><2> ), .B(n1005), .Y(n1782) );
  OAI21X1 U187 ( .A(n1031), .B(n1005), .C(n1781), .Y(n1266) );
  NAND2X1 U188 ( .A(\mem<27><3> ), .B(n1005), .Y(n1781) );
  OAI21X1 U189 ( .A(n1032), .B(n1005), .C(n1780), .Y(n1265) );
  NAND2X1 U190 ( .A(\mem<27><4> ), .B(n1005), .Y(n1780) );
  OAI21X1 U191 ( .A(n1033), .B(n1005), .C(n1779), .Y(n1264) );
  NAND2X1 U192 ( .A(\mem<27><5> ), .B(n1005), .Y(n1779) );
  OAI21X1 U193 ( .A(n1034), .B(n1005), .C(n1778), .Y(n1263) );
  NAND2X1 U194 ( .A(\mem<27><6> ), .B(n1005), .Y(n1778) );
  OAI21X1 U195 ( .A(n1035), .B(n1005), .C(n1777), .Y(n1262) );
  NAND2X1 U196 ( .A(\mem<27><7> ), .B(n1005), .Y(n1777) );
  NAND3X1 U197 ( .A(n973), .B(n1828), .C(n1776), .Y(n1785) );
  OAI21X1 U198 ( .A(n1036), .B(n1004), .C(n1774), .Y(n1261) );
  NAND2X1 U199 ( .A(\mem<26><0> ), .B(n1004), .Y(n1774) );
  OAI21X1 U200 ( .A(n1037), .B(n1003), .C(n1773), .Y(n1260) );
  NAND2X1 U201 ( .A(\mem<26><1> ), .B(n1004), .Y(n1773) );
  OAI21X1 U202 ( .A(n1038), .B(n1003), .C(n1772), .Y(n1259) );
  NAND2X1 U203 ( .A(\mem<26><2> ), .B(n1004), .Y(n1772) );
  OAI21X1 U204 ( .A(n1039), .B(n1003), .C(n1771), .Y(n1258) );
  NAND2X1 U205 ( .A(\mem<26><3> ), .B(n1004), .Y(n1771) );
  OAI21X1 U206 ( .A(n1040), .B(n1003), .C(n1770), .Y(n1257) );
  NAND2X1 U207 ( .A(\mem<26><4> ), .B(n1004), .Y(n1770) );
  OAI21X1 U208 ( .A(n1041), .B(n1003), .C(n1769), .Y(n1256) );
  NAND2X1 U209 ( .A(\mem<26><5> ), .B(n1004), .Y(n1769) );
  OAI21X1 U210 ( .A(n1042), .B(n1003), .C(n1768), .Y(n1255) );
  NAND2X1 U211 ( .A(\mem<26><6> ), .B(n1004), .Y(n1768) );
  OAI21X1 U212 ( .A(n1043), .B(n1003), .C(n1767), .Y(n1254) );
  NAND2X1 U213 ( .A(\mem<26><7> ), .B(n1004), .Y(n1767) );
  NAND3X1 U214 ( .A(n1806), .B(n1828), .C(n1766), .Y(n1775) );
  OAI21X1 U215 ( .A(n1028), .B(n1002), .C(n1764), .Y(n1253) );
  NAND2X1 U216 ( .A(\mem<25><0> ), .B(n1002), .Y(n1764) );
  OAI21X1 U217 ( .A(n1029), .B(n1002), .C(n1763), .Y(n1252) );
  NAND2X1 U218 ( .A(\mem<25><1> ), .B(n1002), .Y(n1763) );
  OAI21X1 U219 ( .A(n1030), .B(n1002), .C(n1762), .Y(n1251) );
  NAND2X1 U220 ( .A(\mem<25><2> ), .B(n1002), .Y(n1762) );
  OAI21X1 U221 ( .A(n1031), .B(n1002), .C(n1761), .Y(n1250) );
  NAND2X1 U222 ( .A(\mem<25><3> ), .B(n1002), .Y(n1761) );
  OAI21X1 U223 ( .A(n1032), .B(n1002), .C(n1760), .Y(n1249) );
  NAND2X1 U224 ( .A(\mem<25><4> ), .B(n1002), .Y(n1760) );
  OAI21X1 U225 ( .A(n1033), .B(n1002), .C(n1759), .Y(n1248) );
  NAND2X1 U226 ( .A(\mem<25><5> ), .B(n1002), .Y(n1759) );
  OAI21X1 U227 ( .A(n1034), .B(n1002), .C(n1758), .Y(n1247) );
  NAND2X1 U228 ( .A(\mem<25><6> ), .B(n1002), .Y(n1758) );
  OAI21X1 U229 ( .A(n1035), .B(n1002), .C(n1757), .Y(n1246) );
  NAND2X1 U230 ( .A(\mem<25><7> ), .B(n1002), .Y(n1757) );
  NAND3X1 U231 ( .A(n973), .B(n1828), .C(n1756), .Y(n1765) );
  OAI21X1 U232 ( .A(n1036), .B(n1001), .C(n1754), .Y(n1245) );
  NAND2X1 U233 ( .A(\mem<24><0> ), .B(n1001), .Y(n1754) );
  OAI21X1 U234 ( .A(n1037), .B(n1000), .C(n1753), .Y(n1244) );
  NAND2X1 U235 ( .A(\mem<24><1> ), .B(n1001), .Y(n1753) );
  OAI21X1 U236 ( .A(n1038), .B(n1000), .C(n1752), .Y(n1243) );
  NAND2X1 U237 ( .A(\mem<24><2> ), .B(n1001), .Y(n1752) );
  OAI21X1 U238 ( .A(n1039), .B(n1000), .C(n1751), .Y(n1242) );
  NAND2X1 U239 ( .A(\mem<24><3> ), .B(n1001), .Y(n1751) );
  OAI21X1 U240 ( .A(n1040), .B(n1000), .C(n1750), .Y(n1241) );
  NAND2X1 U241 ( .A(\mem<24><4> ), .B(n1001), .Y(n1750) );
  OAI21X1 U242 ( .A(n1041), .B(n1000), .C(n1749), .Y(n1240) );
  NAND2X1 U243 ( .A(\mem<24><5> ), .B(n1001), .Y(n1749) );
  OAI21X1 U244 ( .A(n1042), .B(n1000), .C(n1748), .Y(n1239) );
  NAND2X1 U245 ( .A(\mem<24><6> ), .B(n1001), .Y(n1748) );
  OAI21X1 U246 ( .A(n1043), .B(n1000), .C(n1747), .Y(n1238) );
  NAND2X1 U247 ( .A(\mem<24><7> ), .B(n1001), .Y(n1747) );
  NAND3X1 U248 ( .A(n1786), .B(n1828), .C(n1766), .Y(n1755) );
  OAI21X1 U249 ( .A(n1028), .B(n999), .C(n1745), .Y(n1237) );
  NAND2X1 U250 ( .A(\mem<23><0> ), .B(n999), .Y(n1745) );
  OAI21X1 U251 ( .A(n1029), .B(n999), .C(n1744), .Y(n1236) );
  NAND2X1 U252 ( .A(\mem<23><1> ), .B(n999), .Y(n1744) );
  OAI21X1 U253 ( .A(n1030), .B(n999), .C(n1743), .Y(n1235) );
  NAND2X1 U254 ( .A(\mem<23><2> ), .B(n999), .Y(n1743) );
  OAI21X1 U255 ( .A(n1031), .B(n999), .C(n1742), .Y(n1234) );
  NAND2X1 U256 ( .A(\mem<23><3> ), .B(n999), .Y(n1742) );
  OAI21X1 U257 ( .A(n1032), .B(n999), .C(n1741), .Y(n1233) );
  NAND2X1 U258 ( .A(\mem<23><4> ), .B(n999), .Y(n1741) );
  OAI21X1 U259 ( .A(n1033), .B(n999), .C(n1740), .Y(n1232) );
  NAND2X1 U260 ( .A(\mem<23><5> ), .B(n999), .Y(n1740) );
  OAI21X1 U261 ( .A(n1034), .B(n999), .C(n1739), .Y(n1231) );
  NAND2X1 U262 ( .A(\mem<23><6> ), .B(n999), .Y(n1739) );
  OAI21X1 U263 ( .A(n1035), .B(n999), .C(n1738), .Y(n1230) );
  NAND2X1 U264 ( .A(\mem<23><7> ), .B(n999), .Y(n1738) );
  NAND3X1 U265 ( .A(n973), .B(n1828), .C(n1737), .Y(n1746) );
  OAI21X1 U266 ( .A(n1036), .B(n998), .C(n1735), .Y(n1229) );
  NAND2X1 U267 ( .A(\mem<22><0> ), .B(n998), .Y(n1735) );
  OAI21X1 U268 ( .A(n1037), .B(n998), .C(n1734), .Y(n1228) );
  NAND2X1 U269 ( .A(\mem<22><1> ), .B(n998), .Y(n1734) );
  OAI21X1 U270 ( .A(n1038), .B(n998), .C(n1733), .Y(n1227) );
  NAND2X1 U271 ( .A(\mem<22><2> ), .B(n998), .Y(n1733) );
  OAI21X1 U272 ( .A(n1039), .B(n998), .C(n1732), .Y(n1226) );
  NAND2X1 U273 ( .A(\mem<22><3> ), .B(n998), .Y(n1732) );
  OAI21X1 U274 ( .A(n1040), .B(n998), .C(n1731), .Y(n1225) );
  NAND2X1 U275 ( .A(\mem<22><4> ), .B(n998), .Y(n1731) );
  OAI21X1 U276 ( .A(n1041), .B(n998), .C(n1730), .Y(n1224) );
  NAND2X1 U277 ( .A(\mem<22><5> ), .B(n998), .Y(n1730) );
  OAI21X1 U278 ( .A(n1042), .B(n998), .C(n1729), .Y(n1223) );
  NAND2X1 U279 ( .A(\mem<22><6> ), .B(n998), .Y(n1729) );
  OAI21X1 U280 ( .A(n1043), .B(n998), .C(n1728), .Y(n1222) );
  NAND2X1 U281 ( .A(\mem<22><7> ), .B(n998), .Y(n1728) );
  NAND3X1 U282 ( .A(n1806), .B(n1828), .C(n969), .Y(n1736) );
  OAI21X1 U283 ( .A(n1028), .B(n997), .C(n1726), .Y(n1221) );
  NAND2X1 U284 ( .A(\mem<21><0> ), .B(n997), .Y(n1726) );
  OAI21X1 U285 ( .A(n1029), .B(n997), .C(n1725), .Y(n1220) );
  NAND2X1 U286 ( .A(\mem<21><1> ), .B(n997), .Y(n1725) );
  OAI21X1 U287 ( .A(n1030), .B(n997), .C(n1724), .Y(n1219) );
  NAND2X1 U288 ( .A(\mem<21><2> ), .B(n997), .Y(n1724) );
  OAI21X1 U289 ( .A(n1031), .B(n997), .C(n1723), .Y(n1218) );
  NAND2X1 U290 ( .A(\mem<21><3> ), .B(n997), .Y(n1723) );
  OAI21X1 U291 ( .A(n1032), .B(n997), .C(n1722), .Y(n1217) );
  NAND2X1 U292 ( .A(\mem<21><4> ), .B(n997), .Y(n1722) );
  OAI21X1 U293 ( .A(n1033), .B(n997), .C(n1721), .Y(n1216) );
  NAND2X1 U294 ( .A(\mem<21><5> ), .B(n997), .Y(n1721) );
  OAI21X1 U295 ( .A(n1034), .B(n997), .C(n1720), .Y(n1215) );
  NAND2X1 U296 ( .A(\mem<21><6> ), .B(n997), .Y(n1720) );
  OAI21X1 U297 ( .A(n1035), .B(n997), .C(n1719), .Y(n1214) );
  NAND2X1 U298 ( .A(\mem<21><7> ), .B(n997), .Y(n1719) );
  NAND3X1 U299 ( .A(n973), .B(n1828), .C(n1718), .Y(n1727) );
  OAI21X1 U300 ( .A(n1036), .B(n996), .C(n1716), .Y(n1213) );
  NAND2X1 U301 ( .A(\mem<20><0> ), .B(n996), .Y(n1716) );
  OAI21X1 U302 ( .A(n1037), .B(n996), .C(n1715), .Y(n1212) );
  NAND2X1 U303 ( .A(\mem<20><1> ), .B(n996), .Y(n1715) );
  OAI21X1 U304 ( .A(n1038), .B(n996), .C(n1714), .Y(n1211) );
  NAND2X1 U305 ( .A(\mem<20><2> ), .B(n996), .Y(n1714) );
  OAI21X1 U306 ( .A(n1039), .B(n996), .C(n1713), .Y(n1210) );
  NAND2X1 U307 ( .A(\mem<20><3> ), .B(n996), .Y(n1713) );
  OAI21X1 U308 ( .A(n1040), .B(n996), .C(n1712), .Y(n1209) );
  NAND2X1 U309 ( .A(\mem<20><4> ), .B(n996), .Y(n1712) );
  OAI21X1 U310 ( .A(n1041), .B(n996), .C(n1711), .Y(n1208) );
  NAND2X1 U311 ( .A(\mem<20><5> ), .B(n996), .Y(n1711) );
  OAI21X1 U312 ( .A(n1042), .B(n996), .C(n1710), .Y(n1207) );
  NAND2X1 U313 ( .A(\mem<20><6> ), .B(n996), .Y(n1710) );
  OAI21X1 U314 ( .A(n1043), .B(n996), .C(n1709), .Y(n1206) );
  NAND2X1 U315 ( .A(\mem<20><7> ), .B(n996), .Y(n1709) );
  NAND3X1 U316 ( .A(n1786), .B(n1828), .C(n969), .Y(n1717) );
  OAI21X1 U317 ( .A(n1028), .B(n995), .C(n1707), .Y(n1205) );
  NAND2X1 U318 ( .A(\mem<19><0> ), .B(n995), .Y(n1707) );
  OAI21X1 U319 ( .A(n1029), .B(n995), .C(n1706), .Y(n1204) );
  NAND2X1 U320 ( .A(\mem<19><1> ), .B(n995), .Y(n1706) );
  OAI21X1 U321 ( .A(n1030), .B(n995), .C(n1705), .Y(n1203) );
  NAND2X1 U322 ( .A(\mem<19><2> ), .B(n995), .Y(n1705) );
  OAI21X1 U323 ( .A(n1031), .B(n995), .C(n1704), .Y(n1202) );
  NAND2X1 U324 ( .A(\mem<19><3> ), .B(n995), .Y(n1704) );
  OAI21X1 U325 ( .A(n1032), .B(n995), .C(n1703), .Y(n1201) );
  NAND2X1 U326 ( .A(\mem<19><4> ), .B(n995), .Y(n1703) );
  OAI21X1 U327 ( .A(n1033), .B(n995), .C(n1702), .Y(n1200) );
  NAND2X1 U328 ( .A(\mem<19><5> ), .B(n995), .Y(n1702) );
  OAI21X1 U329 ( .A(n1034), .B(n995), .C(n1701), .Y(n1199) );
  NAND2X1 U330 ( .A(\mem<19><6> ), .B(n995), .Y(n1701) );
  OAI21X1 U331 ( .A(n1035), .B(n995), .C(n1700), .Y(n1198) );
  NAND2X1 U332 ( .A(\mem<19><7> ), .B(n995), .Y(n1700) );
  NAND3X1 U333 ( .A(n973), .B(n1828), .C(n1699), .Y(n1708) );
  OAI21X1 U334 ( .A(n1036), .B(n994), .C(n1697), .Y(n1197) );
  NAND2X1 U335 ( .A(\mem<18><0> ), .B(n994), .Y(n1697) );
  OAI21X1 U336 ( .A(n1037), .B(n994), .C(n1696), .Y(n1196) );
  NAND2X1 U337 ( .A(\mem<18><1> ), .B(n994), .Y(n1696) );
  OAI21X1 U338 ( .A(n1038), .B(n994), .C(n1695), .Y(n1195) );
  NAND2X1 U339 ( .A(\mem<18><2> ), .B(n994), .Y(n1695) );
  OAI21X1 U340 ( .A(n1039), .B(n994), .C(n1694), .Y(n1194) );
  NAND2X1 U341 ( .A(\mem<18><3> ), .B(n994), .Y(n1694) );
  OAI21X1 U342 ( .A(n1040), .B(n994), .C(n1693), .Y(n1193) );
  NAND2X1 U343 ( .A(\mem<18><4> ), .B(n994), .Y(n1693) );
  OAI21X1 U344 ( .A(n1041), .B(n994), .C(n1692), .Y(n1192) );
  NAND2X1 U345 ( .A(\mem<18><5> ), .B(n994), .Y(n1692) );
  OAI21X1 U346 ( .A(n1042), .B(n994), .C(n1691), .Y(n1191) );
  NAND2X1 U347 ( .A(\mem<18><6> ), .B(n994), .Y(n1691) );
  OAI21X1 U348 ( .A(n1043), .B(n994), .C(n1690), .Y(n1190) );
  NAND2X1 U349 ( .A(\mem<18><7> ), .B(n994), .Y(n1690) );
  NAND3X1 U350 ( .A(n1806), .B(n1828), .C(n967), .Y(n1698) );
  OAI21X1 U351 ( .A(n1028), .B(n993), .C(n1688), .Y(n1189) );
  NAND2X1 U352 ( .A(\mem<17><0> ), .B(n993), .Y(n1688) );
  OAI21X1 U353 ( .A(n1029), .B(n993), .C(n1687), .Y(n1188) );
  NAND2X1 U354 ( .A(\mem<17><1> ), .B(n993), .Y(n1687) );
  OAI21X1 U355 ( .A(n1030), .B(n993), .C(n1686), .Y(n1187) );
  NAND2X1 U356 ( .A(\mem<17><2> ), .B(n993), .Y(n1686) );
  OAI21X1 U357 ( .A(n1031), .B(n993), .C(n1685), .Y(n1186) );
  NAND2X1 U358 ( .A(\mem<17><3> ), .B(n993), .Y(n1685) );
  OAI21X1 U359 ( .A(n1032), .B(n993), .C(n1684), .Y(n1185) );
  NAND2X1 U360 ( .A(\mem<17><4> ), .B(n993), .Y(n1684) );
  OAI21X1 U361 ( .A(n1033), .B(n993), .C(n1683), .Y(n1184) );
  NAND2X1 U362 ( .A(\mem<17><5> ), .B(n993), .Y(n1683) );
  OAI21X1 U363 ( .A(n1034), .B(n993), .C(n1682), .Y(n1183) );
  NAND2X1 U364 ( .A(\mem<17><6> ), .B(n993), .Y(n1682) );
  OAI21X1 U365 ( .A(n1035), .B(n993), .C(n1681), .Y(n1182) );
  NAND2X1 U366 ( .A(\mem<17><7> ), .B(n993), .Y(n1681) );
  NAND3X1 U367 ( .A(n973), .B(n1828), .C(n1680), .Y(n1689) );
  OAI21X1 U368 ( .A(n1036), .B(n992), .C(n1678), .Y(n1181) );
  NAND2X1 U369 ( .A(\mem<16><0> ), .B(n992), .Y(n1678) );
  OAI21X1 U370 ( .A(n1037), .B(n992), .C(n1677), .Y(n1180) );
  NAND2X1 U371 ( .A(\mem<16><1> ), .B(n992), .Y(n1677) );
  OAI21X1 U372 ( .A(n1038), .B(n992), .C(n1676), .Y(n1179) );
  NAND2X1 U373 ( .A(\mem<16><2> ), .B(n992), .Y(n1676) );
  OAI21X1 U374 ( .A(n1039), .B(n992), .C(n1675), .Y(n1178) );
  NAND2X1 U375 ( .A(\mem<16><3> ), .B(n992), .Y(n1675) );
  OAI21X1 U376 ( .A(n1040), .B(n992), .C(n1674), .Y(n1177) );
  NAND2X1 U377 ( .A(\mem<16><4> ), .B(n992), .Y(n1674) );
  OAI21X1 U378 ( .A(n1041), .B(n992), .C(n1673), .Y(n1176) );
  NAND2X1 U379 ( .A(\mem<16><5> ), .B(n992), .Y(n1673) );
  OAI21X1 U380 ( .A(n1042), .B(n992), .C(n1672), .Y(n1175) );
  NAND2X1 U381 ( .A(\mem<16><6> ), .B(n992), .Y(n1672) );
  OAI21X1 U382 ( .A(n1043), .B(n992), .C(n1671), .Y(n1174) );
  NAND2X1 U383 ( .A(\mem<16><7> ), .B(n992), .Y(n1671) );
  NAND3X1 U384 ( .A(n1786), .B(n1828), .C(n967), .Y(n1679) );
  OAI21X1 U385 ( .A(n1028), .B(n991), .C(n1669), .Y(n1173) );
  NAND2X1 U386 ( .A(\mem<15><0> ), .B(n991), .Y(n1669) );
  OAI21X1 U387 ( .A(n1029), .B(n991), .C(n1668), .Y(n1172) );
  NAND2X1 U388 ( .A(\mem<15><1> ), .B(n991), .Y(n1668) );
  OAI21X1 U389 ( .A(n1030), .B(n991), .C(n1667), .Y(n1171) );
  NAND2X1 U390 ( .A(\mem<15><2> ), .B(n991), .Y(n1667) );
  OAI21X1 U391 ( .A(n1031), .B(n991), .C(n1666), .Y(n1170) );
  NAND2X1 U392 ( .A(\mem<15><3> ), .B(n991), .Y(n1666) );
  OAI21X1 U393 ( .A(n1032), .B(n991), .C(n1665), .Y(n1169) );
  NAND2X1 U394 ( .A(\mem<15><4> ), .B(n991), .Y(n1665) );
  OAI21X1 U395 ( .A(n1033), .B(n991), .C(n1664), .Y(n1168) );
  NAND2X1 U396 ( .A(\mem<15><5> ), .B(n991), .Y(n1664) );
  OAI21X1 U397 ( .A(n1034), .B(n991), .C(n1663), .Y(n1167) );
  NAND2X1 U398 ( .A(\mem<15><6> ), .B(n991), .Y(n1663) );
  OAI21X1 U399 ( .A(n1035), .B(n991), .C(n1662), .Y(n1166) );
  NAND2X1 U400 ( .A(\mem<15><7> ), .B(n991), .Y(n1662) );
  NAND3X1 U401 ( .A(n973), .B(n1828), .C(n1661), .Y(n1670) );
  OAI21X1 U402 ( .A(n1036), .B(n990), .C(n1659), .Y(n1165) );
  NAND2X1 U403 ( .A(\mem<14><0> ), .B(n990), .Y(n1659) );
  OAI21X1 U404 ( .A(n1037), .B(n989), .C(n1658), .Y(n1164) );
  NAND2X1 U405 ( .A(\mem<14><1> ), .B(n990), .Y(n1658) );
  OAI21X1 U406 ( .A(n1038), .B(n989), .C(n1657), .Y(n1163) );
  NAND2X1 U407 ( .A(\mem<14><2> ), .B(n990), .Y(n1657) );
  OAI21X1 U408 ( .A(n1039), .B(n989), .C(n1656), .Y(n1162) );
  NAND2X1 U409 ( .A(\mem<14><3> ), .B(n990), .Y(n1656) );
  OAI21X1 U410 ( .A(n1040), .B(n989), .C(n1655), .Y(n1161) );
  NAND2X1 U411 ( .A(\mem<14><4> ), .B(n990), .Y(n1655) );
  OAI21X1 U412 ( .A(n1041), .B(n989), .C(n1654), .Y(n1160) );
  NAND2X1 U413 ( .A(\mem<14><5> ), .B(n990), .Y(n1654) );
  OAI21X1 U414 ( .A(n1042), .B(n989), .C(n1653), .Y(n1159) );
  NAND2X1 U415 ( .A(\mem<14><6> ), .B(n990), .Y(n1653) );
  OAI21X1 U416 ( .A(n1043), .B(n989), .C(n1652), .Y(n1158) );
  NAND2X1 U417 ( .A(\mem<14><7> ), .B(n990), .Y(n1652) );
  NAND3X1 U418 ( .A(n1807), .B(n1828), .C(n1651), .Y(n1660) );
  OAI21X1 U419 ( .A(n1028), .B(n988), .C(n1649), .Y(n1157) );
  NAND2X1 U420 ( .A(\mem<13><0> ), .B(n988), .Y(n1649) );
  OAI21X1 U421 ( .A(n1029), .B(n988), .C(n1648), .Y(n1156) );
  NAND2X1 U422 ( .A(\mem<13><1> ), .B(n988), .Y(n1648) );
  OAI21X1 U423 ( .A(n1030), .B(n988), .C(n1647), .Y(n1155) );
  NAND2X1 U424 ( .A(\mem<13><2> ), .B(n988), .Y(n1647) );
  OAI21X1 U425 ( .A(n1031), .B(n988), .C(n1646), .Y(n1154) );
  NAND2X1 U426 ( .A(\mem<13><3> ), .B(n988), .Y(n1646) );
  OAI21X1 U427 ( .A(n1032), .B(n988), .C(n1645), .Y(n1153) );
  NAND2X1 U428 ( .A(\mem<13><4> ), .B(n988), .Y(n1645) );
  OAI21X1 U429 ( .A(n1033), .B(n988), .C(n1644), .Y(n1152) );
  NAND2X1 U430 ( .A(\mem<13><5> ), .B(n988), .Y(n1644) );
  OAI21X1 U431 ( .A(n1034), .B(n988), .C(n1643), .Y(n1151) );
  NAND2X1 U432 ( .A(\mem<13><6> ), .B(n988), .Y(n1643) );
  OAI21X1 U433 ( .A(n1035), .B(n988), .C(n1642), .Y(n1150) );
  NAND2X1 U434 ( .A(\mem<13><7> ), .B(n988), .Y(n1642) );
  NAND3X1 U435 ( .A(n973), .B(n1828), .C(n1641), .Y(n1650) );
  OAI21X1 U436 ( .A(n1036), .B(n987), .C(n1639), .Y(n1149) );
  NAND2X1 U437 ( .A(\mem<12><0> ), .B(n987), .Y(n1639) );
  OAI21X1 U438 ( .A(n1037), .B(n986), .C(n1638), .Y(n1148) );
  NAND2X1 U439 ( .A(\mem<12><1> ), .B(n987), .Y(n1638) );
  OAI21X1 U440 ( .A(n1038), .B(n986), .C(n1637), .Y(n1147) );
  NAND2X1 U441 ( .A(\mem<12><2> ), .B(n987), .Y(n1637) );
  OAI21X1 U442 ( .A(n1039), .B(n986), .C(n1636), .Y(n1146) );
  NAND2X1 U443 ( .A(\mem<12><3> ), .B(n987), .Y(n1636) );
  OAI21X1 U444 ( .A(n1040), .B(n986), .C(n1635), .Y(n1145) );
  NAND2X1 U445 ( .A(\mem<12><4> ), .B(n987), .Y(n1635) );
  OAI21X1 U446 ( .A(n1041), .B(n986), .C(n1634), .Y(n1144) );
  NAND2X1 U447 ( .A(\mem<12><5> ), .B(n987), .Y(n1634) );
  OAI21X1 U448 ( .A(n1042), .B(n986), .C(n1633), .Y(n1143) );
  NAND2X1 U449 ( .A(\mem<12><6> ), .B(n987), .Y(n1633) );
  OAI21X1 U450 ( .A(n1043), .B(n986), .C(n1632), .Y(n1142) );
  NAND2X1 U451 ( .A(\mem<12><7> ), .B(n987), .Y(n1632) );
  NAND3X1 U452 ( .A(n1807), .B(n1828), .C(n1631), .Y(n1640) );
  OAI21X1 U453 ( .A(n1028), .B(n985), .C(n1628), .Y(n1141) );
  NAND2X1 U454 ( .A(\mem<11><0> ), .B(n985), .Y(n1628) );
  OAI21X1 U455 ( .A(n1029), .B(n985), .C(n1627), .Y(n1140) );
  NAND2X1 U456 ( .A(\mem<11><1> ), .B(n985), .Y(n1627) );
  OAI21X1 U457 ( .A(n1030), .B(n985), .C(n1626), .Y(n1139) );
  NAND2X1 U458 ( .A(\mem<11><2> ), .B(n985), .Y(n1626) );
  OAI21X1 U459 ( .A(n1031), .B(n985), .C(n1625), .Y(n1138) );
  NAND2X1 U460 ( .A(\mem<11><3> ), .B(n985), .Y(n1625) );
  OAI21X1 U461 ( .A(n1032), .B(n985), .C(n1624), .Y(n1137) );
  NAND2X1 U462 ( .A(\mem<11><4> ), .B(n985), .Y(n1624) );
  OAI21X1 U463 ( .A(n1033), .B(n985), .C(n1623), .Y(n1136) );
  NAND2X1 U464 ( .A(\mem<11><5> ), .B(n985), .Y(n1623) );
  OAI21X1 U465 ( .A(n1034), .B(n985), .C(n1622), .Y(n1135) );
  NAND2X1 U466 ( .A(\mem<11><6> ), .B(n985), .Y(n1622) );
  OAI21X1 U467 ( .A(n1035), .B(n985), .C(n1621), .Y(n1134) );
  NAND2X1 U468 ( .A(\mem<11><7> ), .B(n985), .Y(n1621) );
  NAND3X1 U469 ( .A(n973), .B(n1828), .C(n1620), .Y(n1629) );
  OAI21X1 U470 ( .A(n1036), .B(n984), .C(n1618), .Y(n1133) );
  NAND2X1 U471 ( .A(\mem<10><0> ), .B(n984), .Y(n1618) );
  OAI21X1 U472 ( .A(n1037), .B(n983), .C(n1617), .Y(n1132) );
  NAND2X1 U473 ( .A(\mem<10><1> ), .B(n984), .Y(n1617) );
  OAI21X1 U474 ( .A(n1038), .B(n983), .C(n1616), .Y(n1131) );
  NAND2X1 U475 ( .A(\mem<10><2> ), .B(n984), .Y(n1616) );
  OAI21X1 U476 ( .A(n1039), .B(n983), .C(n1615), .Y(n1130) );
  NAND2X1 U477 ( .A(\mem<10><3> ), .B(n984), .Y(n1615) );
  OAI21X1 U478 ( .A(n1040), .B(n983), .C(n1614), .Y(n1129) );
  NAND2X1 U479 ( .A(\mem<10><4> ), .B(n984), .Y(n1614) );
  OAI21X1 U480 ( .A(n1041), .B(n983), .C(n1613), .Y(n1128) );
  NAND2X1 U481 ( .A(\mem<10><5> ), .B(n984), .Y(n1613) );
  OAI21X1 U482 ( .A(n1042), .B(n983), .C(n1612), .Y(n1127) );
  NAND2X1 U483 ( .A(\mem<10><6> ), .B(n984), .Y(n1612) );
  OAI21X1 U484 ( .A(n1043), .B(n983), .C(n1611), .Y(n1126) );
  NAND2X1 U485 ( .A(\mem<10><7> ), .B(n984), .Y(n1611) );
  NAND3X1 U486 ( .A(n1766), .B(n1828), .C(n1651), .Y(n1619) );
  OAI21X1 U487 ( .A(n1028), .B(n982), .C(n1609), .Y(n1125) );
  NAND2X1 U488 ( .A(\mem<9><0> ), .B(n982), .Y(n1609) );
  OAI21X1 U489 ( .A(n1029), .B(n982), .C(n1608), .Y(n1124) );
  NAND2X1 U490 ( .A(\mem<9><1> ), .B(n982), .Y(n1608) );
  OAI21X1 U491 ( .A(n1030), .B(n982), .C(n1607), .Y(n1123) );
  NAND2X1 U492 ( .A(\mem<9><2> ), .B(n982), .Y(n1607) );
  OAI21X1 U493 ( .A(n1031), .B(n982), .C(n1606), .Y(n1122) );
  NAND2X1 U494 ( .A(\mem<9><3> ), .B(n982), .Y(n1606) );
  OAI21X1 U495 ( .A(n1032), .B(n982), .C(n1605), .Y(n1121) );
  NAND2X1 U496 ( .A(\mem<9><4> ), .B(n982), .Y(n1605) );
  OAI21X1 U497 ( .A(n1033), .B(n982), .C(n1604), .Y(n1120) );
  NAND2X1 U498 ( .A(\mem<9><5> ), .B(n982), .Y(n1604) );
  OAI21X1 U499 ( .A(n1034), .B(n982), .C(n1603), .Y(n1119) );
  NAND2X1 U500 ( .A(\mem<9><6> ), .B(n982), .Y(n1603) );
  OAI21X1 U501 ( .A(n1035), .B(n982), .C(n1602), .Y(n1118) );
  NAND2X1 U502 ( .A(\mem<9><7> ), .B(n982), .Y(n1602) );
  NAND3X1 U503 ( .A(n973), .B(n1828), .C(n1601), .Y(n1610) );
  OAI21X1 U504 ( .A(n1036), .B(n981), .C(n1599), .Y(n1117) );
  NAND2X1 U505 ( .A(\mem<8><0> ), .B(n981), .Y(n1599) );
  OAI21X1 U506 ( .A(n1037), .B(n980), .C(n1598), .Y(n1116) );
  NAND2X1 U507 ( .A(\mem<8><1> ), .B(n981), .Y(n1598) );
  OAI21X1 U508 ( .A(n1038), .B(n980), .C(n1597), .Y(n1115) );
  NAND2X1 U509 ( .A(\mem<8><2> ), .B(n981), .Y(n1597) );
  OAI21X1 U510 ( .A(n1039), .B(n980), .C(n1596), .Y(n1114) );
  NAND2X1 U511 ( .A(\mem<8><3> ), .B(n981), .Y(n1596) );
  OAI21X1 U512 ( .A(n1040), .B(n980), .C(n1595), .Y(n1113) );
  NAND2X1 U513 ( .A(\mem<8><4> ), .B(n981), .Y(n1595) );
  OAI21X1 U514 ( .A(n1041), .B(n980), .C(n1594), .Y(n1112) );
  NAND2X1 U515 ( .A(\mem<8><5> ), .B(n981), .Y(n1594) );
  OAI21X1 U516 ( .A(n1042), .B(n980), .C(n1593), .Y(n1111) );
  NAND2X1 U517 ( .A(\mem<8><6> ), .B(n981), .Y(n1593) );
  OAI21X1 U518 ( .A(n1043), .B(n980), .C(n1592), .Y(n1110) );
  NAND2X1 U519 ( .A(\mem<8><7> ), .B(n981), .Y(n1592) );
  NAND3X1 U520 ( .A(n1766), .B(n1828), .C(n1631), .Y(n1600) );
  OAI21X1 U521 ( .A(n1028), .B(n979), .C(n1589), .Y(n1109) );
  NAND2X1 U522 ( .A(\mem<7><0> ), .B(n979), .Y(n1589) );
  OAI21X1 U523 ( .A(n1029), .B(n979), .C(n1588), .Y(n1108) );
  NAND2X1 U524 ( .A(\mem<7><1> ), .B(n979), .Y(n1588) );
  OAI21X1 U525 ( .A(n1030), .B(n979), .C(n1587), .Y(n1107) );
  NAND2X1 U526 ( .A(\mem<7><2> ), .B(n979), .Y(n1587) );
  OAI21X1 U527 ( .A(n1031), .B(n979), .C(n1586), .Y(n1106) );
  NAND2X1 U528 ( .A(\mem<7><3> ), .B(n979), .Y(n1586) );
  OAI21X1 U529 ( .A(n1032), .B(n979), .C(n1585), .Y(n1105) );
  NAND2X1 U530 ( .A(\mem<7><4> ), .B(n979), .Y(n1585) );
  OAI21X1 U531 ( .A(n1033), .B(n979), .C(n1584), .Y(n1104) );
  NAND2X1 U532 ( .A(\mem<7><5> ), .B(n979), .Y(n1584) );
  OAI21X1 U533 ( .A(n1034), .B(n979), .C(n1583), .Y(n1103) );
  NAND2X1 U534 ( .A(\mem<7><6> ), .B(n979), .Y(n1583) );
  OAI21X1 U535 ( .A(n1035), .B(n979), .C(n1582), .Y(n1102) );
  NAND2X1 U536 ( .A(\mem<7><7> ), .B(n979), .Y(n1582) );
  NAND3X1 U537 ( .A(n973), .B(n1828), .C(n1581), .Y(n1590) );
  OAI21X1 U538 ( .A(n1036), .B(n978), .C(n1579), .Y(n1101) );
  NAND2X1 U539 ( .A(\mem<6><0> ), .B(n978), .Y(n1579) );
  OAI21X1 U540 ( .A(n1037), .B(n978), .C(n1578), .Y(n1100) );
  NAND2X1 U541 ( .A(\mem<6><1> ), .B(n978), .Y(n1578) );
  OAI21X1 U542 ( .A(n1038), .B(n978), .C(n1577), .Y(n1099) );
  NAND2X1 U543 ( .A(\mem<6><2> ), .B(n978), .Y(n1577) );
  OAI21X1 U544 ( .A(n1039), .B(n978), .C(n1576), .Y(n1098) );
  NAND2X1 U545 ( .A(\mem<6><3> ), .B(n978), .Y(n1576) );
  OAI21X1 U546 ( .A(n1040), .B(n978), .C(n1575), .Y(n1097) );
  NAND2X1 U547 ( .A(\mem<6><4> ), .B(n978), .Y(n1575) );
  OAI21X1 U548 ( .A(n1041), .B(n978), .C(n1574), .Y(n1096) );
  NAND2X1 U549 ( .A(\mem<6><5> ), .B(n978), .Y(n1574) );
  OAI21X1 U550 ( .A(n1042), .B(n978), .C(n1573), .Y(n1095) );
  NAND2X1 U551 ( .A(\mem<6><6> ), .B(n978), .Y(n1573) );
  OAI21X1 U552 ( .A(n1043), .B(n978), .C(n1572), .Y(n1094) );
  NAND2X1 U553 ( .A(\mem<6><7> ), .B(n978), .Y(n1572) );
  NAND3X1 U554 ( .A(n969), .B(n1828), .C(n1651), .Y(n1580) );
  OAI21X1 U555 ( .A(n1028), .B(n977), .C(n1570), .Y(n1093) );
  NAND2X1 U556 ( .A(\mem<5><0> ), .B(n977), .Y(n1570) );
  OAI21X1 U557 ( .A(n1029), .B(n977), .C(n1569), .Y(n1092) );
  NAND2X1 U558 ( .A(\mem<5><1> ), .B(n977), .Y(n1569) );
  OAI21X1 U559 ( .A(n1030), .B(n977), .C(n1568), .Y(n1091) );
  NAND2X1 U560 ( .A(\mem<5><2> ), .B(n977), .Y(n1568) );
  OAI21X1 U561 ( .A(n1031), .B(n977), .C(n1567), .Y(n1090) );
  NAND2X1 U562 ( .A(\mem<5><3> ), .B(n977), .Y(n1567) );
  OAI21X1 U563 ( .A(n1032), .B(n977), .C(n1566), .Y(n1089) );
  NAND2X1 U564 ( .A(\mem<5><4> ), .B(n977), .Y(n1566) );
  OAI21X1 U565 ( .A(n1033), .B(n977), .C(n1565), .Y(n1088) );
  NAND2X1 U566 ( .A(\mem<5><5> ), .B(n977), .Y(n1565) );
  OAI21X1 U567 ( .A(n1034), .B(n977), .C(n1564), .Y(n1087) );
  NAND2X1 U568 ( .A(\mem<5><6> ), .B(n977), .Y(n1564) );
  OAI21X1 U569 ( .A(n1035), .B(n977), .C(n1563), .Y(n1086) );
  NAND2X1 U570 ( .A(\mem<5><7> ), .B(n977), .Y(n1563) );
  NAND3X1 U571 ( .A(n973), .B(n1828), .C(n1562), .Y(n1571) );
  OAI21X1 U572 ( .A(n1036), .B(n976), .C(n1560), .Y(n1085) );
  NAND2X1 U573 ( .A(\mem<4><0> ), .B(n976), .Y(n1560) );
  OAI21X1 U574 ( .A(n1037), .B(n976), .C(n1559), .Y(n1084) );
  NAND2X1 U575 ( .A(\mem<4><1> ), .B(n976), .Y(n1559) );
  OAI21X1 U576 ( .A(n1038), .B(n976), .C(n1558), .Y(n1083) );
  NAND2X1 U577 ( .A(\mem<4><2> ), .B(n976), .Y(n1558) );
  OAI21X1 U578 ( .A(n1039), .B(n976), .C(n1557), .Y(n1082) );
  NAND2X1 U579 ( .A(\mem<4><3> ), .B(n976), .Y(n1557) );
  OAI21X1 U580 ( .A(n1040), .B(n976), .C(n1556), .Y(n1081) );
  NAND2X1 U581 ( .A(\mem<4><4> ), .B(n976), .Y(n1556) );
  OAI21X1 U582 ( .A(n1041), .B(n976), .C(n1555), .Y(n1080) );
  NAND2X1 U583 ( .A(\mem<4><5> ), .B(n976), .Y(n1555) );
  OAI21X1 U584 ( .A(n1042), .B(n976), .C(n1554), .Y(n1079) );
  NAND2X1 U585 ( .A(\mem<4><6> ), .B(n976), .Y(n1554) );
  OAI21X1 U586 ( .A(n1043), .B(n976), .C(n1553), .Y(n1078) );
  NAND2X1 U587 ( .A(\mem<4><7> ), .B(n976), .Y(n1553) );
  NAND3X1 U588 ( .A(n969), .B(n1828), .C(n1631), .Y(n1561) );
  OAI21X1 U590 ( .A(n1028), .B(n975), .C(n1550), .Y(n1077) );
  NAND2X1 U591 ( .A(\mem<3><0> ), .B(n975), .Y(n1550) );
  OAI21X1 U592 ( .A(n1029), .B(n975), .C(n1549), .Y(n1076) );
  NAND2X1 U593 ( .A(\mem<3><1> ), .B(n975), .Y(n1549) );
  OAI21X1 U594 ( .A(n1030), .B(n975), .C(n1548), .Y(n1075) );
  NAND2X1 U595 ( .A(\mem<3><2> ), .B(n975), .Y(n1548) );
  OAI21X1 U596 ( .A(n1031), .B(n975), .C(n1547), .Y(n1074) );
  NAND2X1 U597 ( .A(\mem<3><3> ), .B(n975), .Y(n1547) );
  OAI21X1 U598 ( .A(n1032), .B(n975), .C(n1546), .Y(n1073) );
  NAND2X1 U599 ( .A(\mem<3><4> ), .B(n975), .Y(n1546) );
  OAI21X1 U600 ( .A(n1033), .B(n975), .C(n1545), .Y(n1072) );
  NAND2X1 U601 ( .A(\mem<3><5> ), .B(n975), .Y(n1545) );
  OAI21X1 U602 ( .A(n1034), .B(n975), .C(n1544), .Y(n1071) );
  NAND2X1 U603 ( .A(\mem<3><6> ), .B(n975), .Y(n1544) );
  OAI21X1 U604 ( .A(n1035), .B(n975), .C(n1543), .Y(n1070) );
  NAND2X1 U605 ( .A(\mem<3><7> ), .B(n975), .Y(n1543) );
  NAND3X1 U606 ( .A(n973), .B(n1828), .C(n1542), .Y(n1551) );
  OAI21X1 U607 ( .A(n1036), .B(n974), .C(n1540), .Y(n1069) );
  NAND2X1 U608 ( .A(\mem<2><0> ), .B(n974), .Y(n1540) );
  OAI21X1 U609 ( .A(n1037), .B(n974), .C(n1539), .Y(n1068) );
  NAND2X1 U610 ( .A(\mem<2><1> ), .B(n974), .Y(n1539) );
  OAI21X1 U611 ( .A(n1038), .B(n974), .C(n1538), .Y(n1067) );
  NAND2X1 U612 ( .A(\mem<2><2> ), .B(n974), .Y(n1538) );
  OAI21X1 U613 ( .A(n1039), .B(n974), .C(n1537), .Y(n1066) );
  NAND2X1 U614 ( .A(\mem<2><3> ), .B(n974), .Y(n1537) );
  OAI21X1 U615 ( .A(n1040), .B(n974), .C(n1536), .Y(n1065) );
  NAND2X1 U616 ( .A(\mem<2><4> ), .B(n974), .Y(n1536) );
  OAI21X1 U617 ( .A(n1041), .B(n974), .C(n1535), .Y(n1064) );
  NAND2X1 U618 ( .A(\mem<2><5> ), .B(n974), .Y(n1535) );
  OAI21X1 U619 ( .A(n1042), .B(n974), .C(n1534), .Y(n1063) );
  NAND2X1 U620 ( .A(\mem<2><6> ), .B(n974), .Y(n1534) );
  OAI21X1 U621 ( .A(n1043), .B(n974), .C(n1533), .Y(n1062) );
  NAND2X1 U622 ( .A(\mem<2><7> ), .B(n974), .Y(n1533) );
  NAND3X1 U623 ( .A(n967), .B(n1828), .C(n1651), .Y(n1541) );
  OAI21X1 U624 ( .A(n1028), .B(n8), .C(n1532), .Y(n1061) );
  NAND2X1 U625 ( .A(\mem<1><0> ), .B(n8), .Y(n1532) );
  OAI21X1 U626 ( .A(n1029), .B(n8), .C(n1531), .Y(n1060) );
  NAND2X1 U627 ( .A(\mem<1><1> ), .B(n8), .Y(n1531) );
  OAI21X1 U628 ( .A(n1030), .B(n8), .C(n1530), .Y(n1059) );
  NAND2X1 U629 ( .A(\mem<1><2> ), .B(n8), .Y(n1530) );
  OAI21X1 U630 ( .A(n1031), .B(n8), .C(n1529), .Y(n1058) );
  NAND2X1 U631 ( .A(\mem<1><3> ), .B(n8), .Y(n1529) );
  OAI21X1 U632 ( .A(n1032), .B(n8), .C(n1528), .Y(n1057) );
  NAND2X1 U633 ( .A(\mem<1><4> ), .B(n8), .Y(n1528) );
  OAI21X1 U634 ( .A(n1033), .B(n8), .C(n1527), .Y(n1056) );
  NAND2X1 U635 ( .A(\mem<1><5> ), .B(n8), .Y(n1527) );
  OAI21X1 U636 ( .A(n1034), .B(n8), .C(n1526), .Y(n1055) );
  NAND2X1 U637 ( .A(\mem<1><6> ), .B(n8), .Y(n1526) );
  OAI21X1 U638 ( .A(n1035), .B(n8), .C(n1525), .Y(n1054) );
  NAND2X1 U639 ( .A(\mem<1><7> ), .B(n8), .Y(n1525) );
  NOR2X1 U641 ( .A(n965), .B(\addr_1c<4> ), .Y(n1818) );
  OAI21X1 U642 ( .A(n1036), .B(n972), .C(n1522), .Y(n1053) );
  NAND2X1 U643 ( .A(\mem<0><0> ), .B(n972), .Y(n1522) );
  OAI21X1 U644 ( .A(n1037), .B(n972), .C(n1521), .Y(n1052) );
  NAND2X1 U645 ( .A(\mem<0><1> ), .B(n972), .Y(n1521) );
  OAI21X1 U646 ( .A(n1038), .B(n972), .C(n1520), .Y(n1051) );
  NAND2X1 U647 ( .A(\mem<0><2> ), .B(n972), .Y(n1520) );
  OAI21X1 U648 ( .A(n1039), .B(n972), .C(n1519), .Y(n1050) );
  NAND2X1 U649 ( .A(\mem<0><3> ), .B(n972), .Y(n1519) );
  OAI21X1 U650 ( .A(n1040), .B(n972), .C(n1518), .Y(n1049) );
  NAND2X1 U651 ( .A(\mem<0><4> ), .B(n972), .Y(n1518) );
  OAI21X1 U652 ( .A(n1041), .B(n972), .C(n1517), .Y(n1048) );
  NAND2X1 U653 ( .A(\mem<0><5> ), .B(n972), .Y(n1517) );
  OAI21X1 U654 ( .A(n1042), .B(n972), .C(n1516), .Y(n1047) );
  NAND2X1 U655 ( .A(\mem<0><6> ), .B(n972), .Y(n1516) );
  OAI21X1 U656 ( .A(n1043), .B(n972), .C(n1515), .Y(n1046) );
  NAND2X1 U657 ( .A(\mem<0><7> ), .B(n972), .Y(n1515) );
  NAND3X1 U658 ( .A(n967), .B(n1828), .C(n1631), .Y(n1523) );
  NOR3X1 U661 ( .A(n1511), .B(\addr_1c<7> ), .C(\addr_1c<6> ), .Y(n1512) );
  NOR3X1 U662 ( .A(n1510), .B(\addr_1c<11> ), .C(\addr_1c<10> ), .Y(n1513) );
  AOI21X1 U663 ( .A(n461), .B(n1509), .C(n963), .Y(n1838) );
  OAI21X1 U665 ( .A(rd), .B(n1508), .C(wr), .Y(n1509) );
  NAND3X1 U667 ( .A(n1507), .B(n1023), .C(n1506), .Y(n1508) );
  NOR3X1 U668 ( .A(rd1), .B(rd3), .C(rd2), .Y(n1506) );
  NOR2X1 U669 ( .A(wr3), .B(wr2), .Y(n1507) );
  AOI21X1 U670 ( .A(n448), .B(n1504), .C(n1014), .Y(\data_out_1c<9> ) );
  NOR3X1 U671 ( .A(n2), .B(n1503), .C(n4), .Y(n1504) );
  AOI22X1 U673 ( .A(\mem<16><1> ), .B(n1786), .C(\mem<0><1> ), .D(n1631), .Y(
        n1501) );
  AOI22X1 U674 ( .A(\mem<18><1> ), .B(n1806), .C(\mem<2><1> ), .D(n1651), .Y(
        n1502) );
  AOI22X1 U676 ( .A(\mem<20><1> ), .B(n1786), .C(\mem<4><1> ), .D(n1631), .Y(
        n1499) );
  AOI22X1 U677 ( .A(\mem<22><1> ), .B(n1806), .C(\mem<6><1> ), .D(n1651), .Y(
        n1500) );
  AOI22X1 U678 ( .A(n1591), .B(n892), .C(n1630), .D(n932), .Y(n1505) );
  AOI22X1 U680 ( .A(\mem<28><1> ), .B(n1786), .C(\mem<12><1> ), .D(n1631), .Y(
        n1497) );
  AOI22X1 U681 ( .A(\mem<30><1> ), .B(n1806), .C(\mem<14><1> ), .D(n1651), .Y(
        n1498) );
  AOI22X1 U683 ( .A(\mem<24><1> ), .B(n1786), .C(\mem<8><1> ), .D(n1631), .Y(
        n1495) );
  AOI22X1 U684 ( .A(\mem<26><1> ), .B(n1806), .C(\mem<10><1> ), .D(n1651), .Y(
        n1496) );
  AOI21X1 U685 ( .A(n447), .B(n1493), .C(n1014), .Y(\data_out_1c<8> ) );
  NOR3X1 U686 ( .A(n939), .B(n1491), .C(n949), .Y(n1493) );
  AOI21X1 U687 ( .A(n1489), .B(n1488), .C(n971), .Y(n1490) );
  AOI22X1 U688 ( .A(\mem<16><0> ), .B(n1786), .C(\mem<0><0> ), .D(n1631), .Y(
        n1488) );
  AOI22X1 U689 ( .A(\mem<18><0> ), .B(n1806), .C(\mem<2><0> ), .D(n1651), .Y(
        n1489) );
  AOI21X1 U690 ( .A(n1487), .B(n1486), .C(n970), .Y(n1492) );
  AOI22X1 U691 ( .A(\mem<20><0> ), .B(n1786), .C(\mem<4><0> ), .D(n1631), .Y(
        n1486) );
  AOI22X1 U692 ( .A(\mem<22><0> ), .B(n1806), .C(\mem<6><0> ), .D(n1651), .Y(
        n1487) );
  AOI22X1 U693 ( .A(n1591), .B(n890), .C(n1630), .D(n930), .Y(n1494) );
  AOI22X1 U695 ( .A(\mem<28><0> ), .B(n1786), .C(\mem<12><0> ), .D(n1631), .Y(
        n1484) );
  AOI22X1 U696 ( .A(\mem<30><0> ), .B(n1806), .C(\mem<14><0> ), .D(n1651), .Y(
        n1485) );
  AOI22X1 U698 ( .A(\mem<24><0> ), .B(n1786), .C(\mem<8><0> ), .D(n1631), .Y(
        n1482) );
  AOI22X1 U699 ( .A(\mem<26><0> ), .B(n1806), .C(\mem<10><0> ), .D(n1651), .Y(
        n1483) );
  OAI21X1 U700 ( .A(n23), .B(n50), .C(rd1), .Y(n1481) );
  AOI22X1 U702 ( .A(\mem<17><7> ), .B(n1680), .C(\mem<19><7> ), .D(n1699), .Y(
        n1476) );
  AOI22X1 U703 ( .A(\mem<21><7> ), .B(n1718), .C(\mem<23><7> ), .D(n1737), .Y(
        n1477) );
  AOI22X1 U704 ( .A(\mem<25><7> ), .B(n1756), .C(\mem<27><7> ), .D(n1776), .Y(
        n1479) );
  AOI22X1 U705 ( .A(\mem<29><7> ), .B(n1796), .C(\mem<31><7> ), .D(n1817), .Y(
        n1480) );
  AOI22X1 U707 ( .A(\mem<1><7> ), .B(n1524), .C(\mem<3><7> ), .D(n1542), .Y(
        n1471) );
  AOI22X1 U708 ( .A(\mem<5><7> ), .B(n1562), .C(\mem<7><7> ), .D(n1581), .Y(
        n1472) );
  AOI22X1 U709 ( .A(\mem<9><7> ), .B(n1601), .C(\mem<11><7> ), .D(n1620), .Y(
        n1474) );
  AOI22X1 U710 ( .A(\mem<13><7> ), .B(n1641), .C(\mem<15><7> ), .D(n1661), .Y(
        n1475) );
  OAI21X1 U711 ( .A(n21), .B(n37), .C(rd1), .Y(n1470) );
  AOI22X1 U713 ( .A(\mem<17><6> ), .B(n1680), .C(\mem<19><6> ), .D(n1699), .Y(
        n1465) );
  AOI22X1 U714 ( .A(\mem<21><6> ), .B(n1718), .C(\mem<23><6> ), .D(n1737), .Y(
        n1466) );
  AOI22X1 U715 ( .A(\mem<25><6> ), .B(n1756), .C(\mem<27><6> ), .D(n1776), .Y(
        n1468) );
  AOI22X1 U716 ( .A(\mem<29><6> ), .B(n1796), .C(\mem<31><6> ), .D(n1817), .Y(
        n1469) );
  AOI22X1 U718 ( .A(\mem<1><6> ), .B(n1524), .C(\mem<3><6> ), .D(n1542), .Y(
        n1460) );
  AOI22X1 U719 ( .A(\mem<5><6> ), .B(n1562), .C(\mem<7><6> ), .D(n1581), .Y(
        n1461) );
  AOI22X1 U720 ( .A(\mem<9><6> ), .B(n1601), .C(\mem<11><6> ), .D(n1620), .Y(
        n1463) );
  AOI22X1 U721 ( .A(\mem<13><6> ), .B(n1641), .C(\mem<15><6> ), .D(n1661), .Y(
        n1464) );
  OAI21X1 U722 ( .A(n19), .B(n35), .C(rd1), .Y(n1459) );
  AOI22X1 U724 ( .A(\mem<17><5> ), .B(n1680), .C(\mem<19><5> ), .D(n1699), .Y(
        n1454) );
  AOI22X1 U725 ( .A(\mem<21><5> ), .B(n1718), .C(\mem<23><5> ), .D(n1737), .Y(
        n1455) );
  AOI22X1 U726 ( .A(\mem<25><5> ), .B(n1756), .C(\mem<27><5> ), .D(n1776), .Y(
        n1457) );
  AOI22X1 U727 ( .A(\mem<29><5> ), .B(n1796), .C(\mem<31><5> ), .D(n1817), .Y(
        n1458) );
  AOI22X1 U729 ( .A(\mem<1><5> ), .B(n1524), .C(\mem<3><5> ), .D(n1542), .Y(
        n1449) );
  AOI22X1 U730 ( .A(\mem<5><5> ), .B(n1562), .C(\mem<7><5> ), .D(n1581), .Y(
        n1450) );
  AOI22X1 U731 ( .A(\mem<9><5> ), .B(n1601), .C(\mem<11><5> ), .D(n1620), .Y(
        n1452) );
  AOI22X1 U732 ( .A(\mem<13><5> ), .B(n1641), .C(\mem<15><5> ), .D(n1661), .Y(
        n1453) );
  OAI21X1 U733 ( .A(n17), .B(n33), .C(rd1), .Y(n1448) );
  AOI22X1 U735 ( .A(\mem<17><4> ), .B(n1680), .C(\mem<19><4> ), .D(n1699), .Y(
        n1443) );
  AOI22X1 U736 ( .A(\mem<21><4> ), .B(n1718), .C(\mem<23><4> ), .D(n1737), .Y(
        n1444) );
  AOI22X1 U737 ( .A(\mem<25><4> ), .B(n1756), .C(\mem<27><4> ), .D(n1776), .Y(
        n1446) );
  AOI22X1 U738 ( .A(\mem<29><4> ), .B(n1796), .C(\mem<31><4> ), .D(n1817), .Y(
        n1447) );
  AOI22X1 U740 ( .A(\mem<1><4> ), .B(n1524), .C(\mem<3><4> ), .D(n1542), .Y(
        n1438) );
  AOI22X1 U741 ( .A(\mem<5><4> ), .B(n1562), .C(\mem<7><4> ), .D(n1581), .Y(
        n1439) );
  AOI22X1 U742 ( .A(\mem<9><4> ), .B(n1601), .C(\mem<11><4> ), .D(n1620), .Y(
        n1441) );
  AOI22X1 U743 ( .A(\mem<13><4> ), .B(n1641), .C(\mem<15><4> ), .D(n1661), .Y(
        n1442) );
  OAI21X1 U744 ( .A(n15), .B(n31), .C(rd1), .Y(n1437) );
  AOI22X1 U746 ( .A(\mem<17><3> ), .B(n1680), .C(\mem<19><3> ), .D(n1699), .Y(
        n1432) );
  AOI22X1 U747 ( .A(\mem<21><3> ), .B(n1718), .C(\mem<23><3> ), .D(n1737), .Y(
        n1433) );
  AOI22X1 U748 ( .A(\mem<25><3> ), .B(n1756), .C(\mem<27><3> ), .D(n1776), .Y(
        n1435) );
  AOI22X1 U749 ( .A(\mem<29><3> ), .B(n1796), .C(\mem<31><3> ), .D(n1817), .Y(
        n1436) );
  AOI22X1 U751 ( .A(\mem<1><3> ), .B(n1524), .C(\mem<3><3> ), .D(n1542), .Y(
        n1427) );
  AOI22X1 U752 ( .A(\mem<5><3> ), .B(n1562), .C(\mem<7><3> ), .D(n1581), .Y(
        n1428) );
  AOI22X1 U753 ( .A(\mem<9><3> ), .B(n1601), .C(\mem<11><3> ), .D(n1620), .Y(
        n1430) );
  AOI22X1 U754 ( .A(\mem<13><3> ), .B(n1641), .C(\mem<15><3> ), .D(n1661), .Y(
        n1431) );
  OAI21X1 U755 ( .A(n13), .B(n29), .C(rd1), .Y(n1426) );
  AOI22X1 U757 ( .A(\mem<17><2> ), .B(n1680), .C(\mem<19><2> ), .D(n1699), .Y(
        n1421) );
  AOI22X1 U758 ( .A(\mem<21><2> ), .B(n1718), .C(\mem<23><2> ), .D(n1737), .Y(
        n1422) );
  AOI22X1 U759 ( .A(\mem<25><2> ), .B(n1756), .C(\mem<27><2> ), .D(n1776), .Y(
        n1424) );
  AOI22X1 U760 ( .A(\mem<29><2> ), .B(n1796), .C(\mem<31><2> ), .D(n1817), .Y(
        n1425) );
  AOI22X1 U762 ( .A(\mem<1><2> ), .B(n1524), .C(\mem<3><2> ), .D(n1542), .Y(
        n1416) );
  AOI22X1 U763 ( .A(\mem<5><2> ), .B(n1562), .C(\mem<7><2> ), .D(n1581), .Y(
        n1417) );
  AOI22X1 U764 ( .A(\mem<9><2> ), .B(n1601), .C(\mem<11><2> ), .D(n1620), .Y(
        n1419) );
  AOI22X1 U765 ( .A(\mem<13><2> ), .B(n1641), .C(\mem<15><2> ), .D(n1661), .Y(
        n1420) );
  OAI21X1 U766 ( .A(n11), .B(n27), .C(rd1), .Y(n1415) );
  AOI22X1 U768 ( .A(\mem<17><1> ), .B(n1680), .C(\mem<19><1> ), .D(n1699), .Y(
        n1410) );
  AOI22X1 U769 ( .A(\mem<21><1> ), .B(n1718), .C(\mem<23><1> ), .D(n1737), .Y(
        n1411) );
  AOI22X1 U770 ( .A(\mem<25><1> ), .B(n1756), .C(\mem<27><1> ), .D(n1776), .Y(
        n1413) );
  AOI22X1 U771 ( .A(\mem<29><1> ), .B(n1796), .C(\mem<31><1> ), .D(n1817), .Y(
        n1414) );
  AOI22X1 U773 ( .A(\mem<1><1> ), .B(n1524), .C(\mem<3><1> ), .D(n1542), .Y(
        n1405) );
  AOI22X1 U774 ( .A(\mem<5><1> ), .B(n1562), .C(\mem<7><1> ), .D(n1581), .Y(
        n1406) );
  AOI22X1 U775 ( .A(\mem<9><1> ), .B(n1601), .C(\mem<11><1> ), .D(n1620), .Y(
        n1408) );
  AOI22X1 U776 ( .A(\mem<13><1> ), .B(n1641), .C(\mem<15><1> ), .D(n1661), .Y(
        n1409) );
  AOI21X1 U777 ( .A(n435), .B(n1403), .C(n1014), .Y(\data_out_1c<15> ) );
  NOR3X1 U778 ( .A(n938), .B(n1401), .C(n948), .Y(n1403) );
  AOI21X1 U779 ( .A(n1399), .B(n1398), .C(n971), .Y(n1400) );
  AOI22X1 U780 ( .A(\mem<16><7> ), .B(n1786), .C(\mem<0><7> ), .D(n1631), .Y(
        n1398) );
  AOI22X1 U781 ( .A(\mem<18><7> ), .B(n1806), .C(\mem<2><7> ), .D(n1651), .Y(
        n1399) );
  AOI21X1 U782 ( .A(n1397), .B(n1396), .C(n970), .Y(n1402) );
  AOI22X1 U783 ( .A(\mem<20><7> ), .B(n1786), .C(\mem<4><7> ), .D(n1631), .Y(
        n1396) );
  AOI22X1 U784 ( .A(\mem<22><7> ), .B(n1806), .C(\mem<6><7> ), .D(n1651), .Y(
        n1397) );
  AOI22X1 U785 ( .A(n1591), .B(n888), .C(n1630), .D(n928), .Y(n1404) );
  AOI22X1 U787 ( .A(\mem<28><7> ), .B(n1786), .C(\mem<12><7> ), .D(n1631), .Y(
        n1394) );
  AOI22X1 U788 ( .A(\mem<30><7> ), .B(n1806), .C(\mem<14><7> ), .D(n1651), .Y(
        n1395) );
  AOI22X1 U790 ( .A(\mem<24><7> ), .B(n1786), .C(\mem<8><7> ), .D(n1631), .Y(
        n1392) );
  AOI22X1 U791 ( .A(\mem<26><7> ), .B(n1806), .C(\mem<10><7> ), .D(n1651), .Y(
        n1393) );
  AOI21X1 U792 ( .A(n434), .B(n1390), .C(n1014), .Y(\data_out_1c<14> ) );
  NOR3X1 U793 ( .A(n937), .B(n1388), .C(n947), .Y(n1390) );
  AOI21X1 U794 ( .A(n1386), .B(n1385), .C(n971), .Y(n1387) );
  AOI22X1 U795 ( .A(\mem<16><6> ), .B(n1786), .C(\mem<0><6> ), .D(n1631), .Y(
        n1385) );
  AOI22X1 U796 ( .A(\mem<18><6> ), .B(n1806), .C(\mem<2><6> ), .D(n1651), .Y(
        n1386) );
  AOI21X1 U797 ( .A(n1384), .B(n1383), .C(n970), .Y(n1389) );
  AOI22X1 U798 ( .A(\mem<20><6> ), .B(n1786), .C(\mem<4><6> ), .D(n1631), .Y(
        n1383) );
  AOI22X1 U799 ( .A(\mem<22><6> ), .B(n1806), .C(\mem<6><6> ), .D(n1651), .Y(
        n1384) );
  AOI22X1 U800 ( .A(n1591), .B(n886), .C(n1630), .D(n926), .Y(n1391) );
  AOI22X1 U802 ( .A(\mem<28><6> ), .B(n1786), .C(\mem<12><6> ), .D(n1631), .Y(
        n1381) );
  AOI22X1 U803 ( .A(\mem<30><6> ), .B(n1806), .C(\mem<14><6> ), .D(n1651), .Y(
        n1382) );
  AOI22X1 U805 ( .A(\mem<24><6> ), .B(n1786), .C(\mem<8><6> ), .D(n1631), .Y(
        n1379) );
  AOI22X1 U806 ( .A(\mem<26><6> ), .B(n1806), .C(\mem<10><6> ), .D(n1651), .Y(
        n1380) );
  AOI21X1 U807 ( .A(n422), .B(n1377), .C(n1014), .Y(\data_out_1c<13> ) );
  NOR3X1 U808 ( .A(n936), .B(n1375), .C(n946), .Y(n1377) );
  AOI21X1 U809 ( .A(n1373), .B(n1372), .C(n971), .Y(n1374) );
  AOI22X1 U810 ( .A(\mem<16><5> ), .B(n1786), .C(\mem<0><5> ), .D(n1631), .Y(
        n1372) );
  AOI22X1 U811 ( .A(\mem<18><5> ), .B(n1806), .C(\mem<2><5> ), .D(n1651), .Y(
        n1373) );
  AOI21X1 U812 ( .A(n1371), .B(n1370), .C(n970), .Y(n1376) );
  AOI22X1 U813 ( .A(\mem<20><5> ), .B(n1786), .C(\mem<4><5> ), .D(n1631), .Y(
        n1370) );
  AOI22X1 U814 ( .A(\mem<22><5> ), .B(n1806), .C(\mem<6><5> ), .D(n1651), .Y(
        n1371) );
  AOI22X1 U815 ( .A(n1591), .B(n884), .C(n1630), .D(n924), .Y(n1378) );
  AOI22X1 U817 ( .A(\mem<28><5> ), .B(n1786), .C(\mem<12><5> ), .D(n1631), .Y(
        n1368) );
  AOI22X1 U818 ( .A(\mem<30><5> ), .B(n1806), .C(\mem<14><5> ), .D(n1651), .Y(
        n1369) );
  AOI22X1 U820 ( .A(\mem<24><5> ), .B(n1786), .C(\mem<8><5> ), .D(n1631), .Y(
        n1366) );
  AOI22X1 U821 ( .A(\mem<26><5> ), .B(n1806), .C(\mem<10><5> ), .D(n1651), .Y(
        n1367) );
  AOI21X1 U822 ( .A(n421), .B(n1364), .C(n1014), .Y(\data_out_1c<12> ) );
  NOR3X1 U823 ( .A(n935), .B(n1362), .C(n945), .Y(n1364) );
  AOI21X1 U824 ( .A(n1360), .B(n1359), .C(n971), .Y(n1361) );
  AOI22X1 U825 ( .A(\mem<16><4> ), .B(n1786), .C(\mem<0><4> ), .D(n1631), .Y(
        n1359) );
  AOI22X1 U826 ( .A(\mem<18><4> ), .B(n1806), .C(\mem<2><4> ), .D(n1651), .Y(
        n1360) );
  AOI21X1 U827 ( .A(n1358), .B(n1357), .C(n970), .Y(n1363) );
  AOI22X1 U828 ( .A(\mem<20><4> ), .B(n1786), .C(\mem<4><4> ), .D(n1631), .Y(
        n1357) );
  AOI22X1 U829 ( .A(\mem<22><4> ), .B(n1806), .C(\mem<6><4> ), .D(n1651), .Y(
        n1358) );
  AOI22X1 U830 ( .A(n1591), .B(n882), .C(n1630), .D(n922), .Y(n1365) );
  AOI22X1 U832 ( .A(\mem<28><4> ), .B(n1786), .C(\mem<12><4> ), .D(n1631), .Y(
        n1355) );
  AOI22X1 U833 ( .A(\mem<30><4> ), .B(n1806), .C(\mem<14><4> ), .D(n1651), .Y(
        n1356) );
  AOI22X1 U835 ( .A(\mem<24><4> ), .B(n1786), .C(\mem<8><4> ), .D(n1631), .Y(
        n1353) );
  AOI22X1 U836 ( .A(\mem<26><4> ), .B(n1806), .C(\mem<10><4> ), .D(n1651), .Y(
        n1354) );
  AOI21X1 U837 ( .A(n409), .B(n1351), .C(n1014), .Y(\data_out_1c<11> ) );
  NOR3X1 U838 ( .A(n934), .B(n1349), .C(n944), .Y(n1351) );
  AOI21X1 U839 ( .A(n1347), .B(n1346), .C(n971), .Y(n1348) );
  AOI22X1 U840 ( .A(\mem<16><3> ), .B(n1786), .C(\mem<0><3> ), .D(n1631), .Y(
        n1346) );
  AOI22X1 U841 ( .A(\mem<18><3> ), .B(n1806), .C(\mem<2><3> ), .D(n1651), .Y(
        n1347) );
  AOI21X1 U842 ( .A(n1345), .B(n1344), .C(n970), .Y(n1350) );
  AOI22X1 U843 ( .A(\mem<20><3> ), .B(n1786), .C(\mem<4><3> ), .D(n1631), .Y(
        n1344) );
  AOI22X1 U844 ( .A(\mem<22><3> ), .B(n1806), .C(\mem<6><3> ), .D(n1651), .Y(
        n1345) );
  AOI22X1 U845 ( .A(n1591), .B(n880), .C(n1630), .D(n920), .Y(n1352) );
  AOI22X1 U847 ( .A(\mem<28><3> ), .B(n1786), .C(\mem<12><3> ), .D(n1631), .Y(
        n1342) );
  AOI22X1 U848 ( .A(\mem<30><3> ), .B(n1806), .C(\mem<14><3> ), .D(n1651), .Y(
        n1343) );
  AOI22X1 U850 ( .A(\mem<24><3> ), .B(n1786), .C(\mem<8><3> ), .D(n1631), .Y(
        n1340) );
  AOI22X1 U851 ( .A(\mem<26><3> ), .B(n1806), .C(\mem<10><3> ), .D(n1651), .Y(
        n1341) );
  AOI21X1 U852 ( .A(n408), .B(n1338), .C(n1014), .Y(\data_out_1c<10> ) );
  NOR3X1 U853 ( .A(n933), .B(n1336), .C(n943), .Y(n1338) );
  AOI21X1 U854 ( .A(n1334), .B(n1333), .C(n971), .Y(n1335) );
  AOI22X1 U855 ( .A(\mem<16><2> ), .B(n1786), .C(\mem<0><2> ), .D(n1631), .Y(
        n1333) );
  AOI22X1 U856 ( .A(\mem<18><2> ), .B(n1806), .C(\mem<2><2> ), .D(n1651), .Y(
        n1334) );
  AOI21X1 U857 ( .A(n1332), .B(n1331), .C(n970), .Y(n1337) );
  AOI22X1 U858 ( .A(\mem<20><2> ), .B(n1786), .C(\mem<4><2> ), .D(n1631), .Y(
        n1331) );
  AOI22X1 U859 ( .A(\mem<22><2> ), .B(n1806), .C(\mem<6><2> ), .D(n1651), .Y(
        n1332) );
  AOI22X1 U860 ( .A(n1591), .B(n878), .C(n1630), .D(n918), .Y(n1339) );
  AOI22X1 U862 ( .A(\mem<28><2> ), .B(n1786), .C(\mem<12><2> ), .D(n1631), .Y(
        n1329) );
  AOI22X1 U863 ( .A(\mem<30><2> ), .B(n1806), .C(\mem<14><2> ), .D(n1651), .Y(
        n1330) );
  AOI22X1 U865 ( .A(\mem<24><2> ), .B(n1786), .C(\mem<8><2> ), .D(n1631), .Y(
        n1327) );
  AOI22X1 U866 ( .A(\mem<26><2> ), .B(n1806), .C(\mem<10><2> ), .D(n1651), .Y(
        n1328) );
  NOR2X1 U867 ( .A(\addr_1c<3> ), .B(\addr_1c<4> ), .Y(n1326) );
  NOR2X1 U868 ( .A(n1027), .B(\addr_1c<4> ), .Y(n1325) );
  OAI21X1 U869 ( .A(n9), .B(n25), .C(rd1), .Y(n1324) );
  AOI22X1 U871 ( .A(\mem<17><0> ), .B(n1680), .C(\mem<19><0> ), .D(n1699), .Y(
        n1319) );
  AOI22X1 U872 ( .A(\mem<21><0> ), .B(n1718), .C(\mem<23><0> ), .D(n1737), .Y(
        n1320) );
  AOI22X1 U873 ( .A(\mem<25><0> ), .B(n1756), .C(\mem<27><0> ), .D(n1776), .Y(
        n1322) );
  AOI22X1 U874 ( .A(\mem<29><0> ), .B(n1796), .C(\mem<31><0> ), .D(n1817), .Y(
        n1323) );
  AOI22X1 U876 ( .A(\mem<1><0> ), .B(n1524), .C(\mem<3><0> ), .D(n1542), .Y(
        n1312) );
  NAND2X1 U877 ( .A(n1025), .B(n1026), .Y(n1514) );
  AOI22X1 U878 ( .A(\mem<5><0> ), .B(n1562), .C(\mem<7><0> ), .D(n1581), .Y(
        n1313) );
  NAND2X1 U879 ( .A(\addr_1c<1> ), .B(n1026), .Y(n1552) );
  AOI22X1 U880 ( .A(\mem<9><0> ), .B(n1601), .C(\mem<11><0> ), .D(n1620), .Y(
        n1315) );
  AOI22X1 U881 ( .A(\mem<13><0> ), .B(n1641), .C(\mem<15><0> ), .D(n1661), .Y(
        n1316) );
  dff_105 ff0 ( .q(rd1), .d(rd0), .clk(clk), .rst(n1012) );
  dff_104 ff1 ( .q(wr1), .d(wr0), .clk(clk), .rst(n1012) );
  dff_103 \reg0[0]  ( .q(\addr_1c<0> ), .d(\addr<0> ), .clk(clk), .rst(n1012)
         );
  dff_102 \reg0[1]  ( .q(\addr_1c<1> ), .d(\addr<1> ), .clk(clk), .rst(n1012)
         );
  dff_101 \reg0[2]  ( .q(\addr_1c<2> ), .d(\addr<2> ), .clk(clk), .rst(n1012)
         );
  dff_100 \reg0[3]  ( .q(\addr_1c<3> ), .d(\addr<3> ), .clk(clk), .rst(n1012)
         );
  dff_99 \reg0[4]  ( .q(\addr_1c<4> ), .d(\addr<4> ), .clk(clk), .rst(n1012)
         );
  dff_98 \reg0[5]  ( .q(\addr_1c<5> ), .d(\addr<5> ), .clk(clk), .rst(n1012)
         );
  dff_97 \reg0[6]  ( .q(\addr_1c<6> ), .d(\addr<6> ), .clk(clk), .rst(n1012)
         );
  dff_96 \reg0[7]  ( .q(\addr_1c<7> ), .d(\addr<7> ), .clk(clk), .rst(n1012)
         );
  dff_95 \reg0[8]  ( .q(\addr_1c<8> ), .d(\addr<8> ), .clk(clk), .rst(n1012)
         );
  dff_94 \reg0[9]  ( .q(\addr_1c<9> ), .d(\addr<9> ), .clk(clk), .rst(n1012)
         );
  dff_93 \reg0[10]  ( .q(\addr_1c<10> ), .d(\addr<10> ), .clk(clk), .rst(n1012) );
  dff_92 \reg0[11]  ( .q(\addr_1c<11> ), .d(\addr<11> ), .clk(clk), .rst(n1012) );
  dff_91 \reg0[12]  ( .q(\addr_1c<12> ), .d(\addr<12> ), .clk(clk), .rst(n1012) );
  dff_90 \reg1[0]  ( .q(\data_in_1c<0> ), .d(\data_in<0> ), .clk(clk), .rst(
        n1012) );
  dff_89 \reg1[1]  ( .q(\data_in_1c<1> ), .d(\data_in<1> ), .clk(clk), .rst(
        n1012) );
  dff_88 \reg1[2]  ( .q(\data_in_1c<2> ), .d(\data_in<2> ), .clk(clk), .rst(
        n1012) );
  dff_87 \reg1[3]  ( .q(\data_in_1c<3> ), .d(\data_in<3> ), .clk(clk), .rst(
        n1012) );
  dff_86 \reg1[4]  ( .q(\data_in_1c<4> ), .d(\data_in<4> ), .clk(clk), .rst(
        n1012) );
  dff_85 \reg1[5]  ( .q(\data_in_1c<5> ), .d(\data_in<5> ), .clk(clk), .rst(
        n1012) );
  dff_84 \reg1[6]  ( .q(\data_in_1c<6> ), .d(\data_in<6> ), .clk(clk), .rst(
        n1012) );
  dff_83 \reg1[7]  ( .q(\data_in_1c<7> ), .d(\data_in<7> ), .clk(clk), .rst(
        n1012) );
  dff_82 \reg1[8]  ( .q(\data_in_1c<8> ), .d(\data_in<8> ), .clk(clk), .rst(
        n1012) );
  dff_81 \reg1[9]  ( .q(\data_in_1c<9> ), .d(\data_in<9> ), .clk(clk), .rst(
        n1012) );
  dff_80 \reg1[10]  ( .q(\data_in_1c<10> ), .d(\data_in<10> ), .clk(clk), 
        .rst(n1012) );
  dff_79 \reg1[11]  ( .q(\data_in_1c<11> ), .d(\data_in<11> ), .clk(clk), 
        .rst(n1012) );
  dff_78 \reg1[12]  ( .q(\data_in_1c<12> ), .d(\data_in<12> ), .clk(clk), 
        .rst(n1012) );
  dff_77 \reg1[13]  ( .q(\data_in_1c<13> ), .d(\data_in<13> ), .clk(clk), 
        .rst(n1012) );
  dff_76 \reg1[14]  ( .q(\data_in_1c<14> ), .d(\data_in<14> ), .clk(clk), 
        .rst(n1012) );
  dff_75 \reg1[15]  ( .q(\data_in_1c<15> ), .d(\data_in<15> ), .clk(clk), 
        .rst(n1012) );
  dff_74 \reg2[0]  ( .q(\data_out<0> ), .d(n1022), .clk(clk), .rst(n1012) );
  dff_73 \reg2[1]  ( .q(\data_out<1> ), .d(n1021), .clk(clk), .rst(n1012) );
  dff_72 \reg2[2]  ( .q(\data_out<2> ), .d(n1020), .clk(clk), .rst(n1012) );
  dff_71 \reg2[3]  ( .q(\data_out<3> ), .d(n1019), .clk(clk), .rst(n1012) );
  dff_70 \reg2[4]  ( .q(\data_out<4> ), .d(n1018), .clk(clk), .rst(n1012) );
  dff_69 \reg2[5]  ( .q(\data_out<5> ), .d(n1017), .clk(clk), .rst(n1012) );
  dff_68 \reg2[6]  ( .q(\data_out<6> ), .d(n1016), .clk(clk), .rst(n1012) );
  dff_67 \reg2[7]  ( .q(\data_out<7> ), .d(n1015), .clk(clk), .rst(n1012) );
  dff_66 \reg2[8]  ( .q(\data_out<8> ), .d(\data_out_1c<8> ), .clk(clk), .rst(
        n1012) );
  dff_65 \reg2[9]  ( .q(\data_out<9> ), .d(\data_out_1c<9> ), .clk(clk), .rst(
        n1012) );
  dff_64 \reg2[10]  ( .q(\data_out<10> ), .d(\data_out_1c<10> ), .clk(clk), 
        .rst(n1012) );
  dff_63 \reg2[11]  ( .q(\data_out<11> ), .d(\data_out_1c<11> ), .clk(clk), 
        .rst(n1012) );
  dff_62 \reg2[12]  ( .q(\data_out<12> ), .d(\data_out_1c<12> ), .clk(clk), 
        .rst(n1012) );
  dff_61 \reg2[13]  ( .q(\data_out<13> ), .d(\data_out_1c<13> ), .clk(clk), 
        .rst(n1012) );
  dff_60 \reg2[14]  ( .q(\data_out<14> ), .d(\data_out_1c<14> ), .clk(clk), 
        .rst(n1012) );
  dff_59 \reg2[15]  ( .q(\data_out<15> ), .d(\data_out_1c<15> ), .clk(clk), 
        .rst(n1012) );
  dff_58 ff2 ( .q(rd2), .d(rd1), .clk(clk), .rst(n1012) );
  dff_57 ff3 ( .q(wr2), .d(wr1), .clk(clk), .rst(n1012) );
  dff_56 ff4 ( .q(rd3), .d(rd2), .clk(clk), .rst(n1012) );
  dff_55 ff5 ( .q(wr3), .d(wr2), .clk(clk), .rst(n1012) );
  INVX1 U2 ( .A(rd), .Y(n1045) );
  OR2X1 U3 ( .A(\addr_1c<5> ), .B(\addr_1c<12> ), .Y(n1510) );
  AND2X1 U4 ( .A(\addr_1c<4> ), .B(n1524), .Y(n1827) );
  INVX1 U5 ( .A(\addr_1c<3> ), .Y(n1027) );
  INVX1 U6 ( .A(\addr_1c<2> ), .Y(n1026) );
  INVX1 U7 ( .A(wr1), .Y(n1023) );
  INVX1 U8 ( .A(\addr_1c<1> ), .Y(n1025) );
  OR2X1 U23 ( .A(\addr_1c<9> ), .B(\addr_1c<8> ), .Y(n1511) );
  AND2X1 U24 ( .A(\addr_1c<3> ), .B(\addr_1c<0> ), .Y(n1318) );
  AND2X1 U25 ( .A(\addr_1c<3> ), .B(n1024), .Y(n1317) );
  AND2X1 U26 ( .A(n1630), .B(n964), .Y(n1807) );
  AND2X1 U27 ( .A(n1591), .B(n964), .Y(n1766) );
  AND2X1 U28 ( .A(\addr_1c<0> ), .B(n1027), .Y(n1311) );
  AND2X1 U29 ( .A(n1024), .B(n1027), .Y(n1310) );
  INVX1 U35 ( .A(\addr_1c<0> ), .Y(n1024) );
  AND2X1 U36 ( .A(\addr_1c<2> ), .B(n1025), .Y(n1591) );
  AND2X1 U37 ( .A(\addr_1c<2> ), .B(\addr_1c<1> ), .Y(n1630) );
  AND2X1 U38 ( .A(n1317), .B(n1630), .Y(n1796) );
  AND2X1 U39 ( .A(n1591), .B(n1318), .Y(n1776) );
  AND2X1 U40 ( .A(n1591), .B(n1317), .Y(n1756) );
  AND2X1 U41 ( .A(n940), .B(n1318), .Y(n1737) );
  AND2X1 U42 ( .A(n940), .B(n1317), .Y(n1718) );
  AND2X1 U43 ( .A(n1318), .B(n950), .Y(n1699) );
  AND2X1 U44 ( .A(n1317), .B(n950), .Y(n1680) );
  AND2X1 U46 ( .A(n1311), .B(n1630), .Y(n1661) );
  AND2X1 U47 ( .A(n1630), .B(n1310), .Y(n1641) );
  AND2X1 U48 ( .A(n1311), .B(n1591), .Y(n1620) );
  AND2X1 U49 ( .A(n1591), .B(n1310), .Y(n1601) );
  AND2X1 U50 ( .A(n1311), .B(n940), .Y(n1581) );
  AND2X1 U51 ( .A(n940), .B(n1310), .Y(n1562) );
  OR2X1 U52 ( .A(n970), .B(n965), .Y(n968) );
  AND2X1 U53 ( .A(n1311), .B(n950), .Y(n1542) );
  OR2X1 U54 ( .A(n965), .B(n971), .Y(n966) );
  AND2X1 U55 ( .A(n1827), .B(\mem<32><0> ), .Y(n1491) );
  AND2X1 U56 ( .A(n1827), .B(\mem<32><1> ), .Y(n1503) );
  AND2X1 U57 ( .A(n1827), .B(\mem<32><2> ), .Y(n1336) );
  AND2X1 U58 ( .A(n1827), .B(\mem<32><3> ), .Y(n1349) );
  AND2X1 U59 ( .A(n1827), .B(\mem<32><4> ), .Y(n1362) );
  AND2X1 U60 ( .A(n1827), .B(\mem<32><5> ), .Y(n1375) );
  AND2X1 U61 ( .A(n1827), .B(\mem<32><6> ), .Y(n1388) );
  AND2X1 U62 ( .A(n1827), .B(\mem<32><7> ), .Y(n1401) );
  INVX1 U63 ( .A(rd1), .Y(n1014) );
  BUFX2 U64 ( .A(n961), .Y(n1010) );
  BUFX2 U65 ( .A(n961), .Y(n1009) );
  BUFX2 U66 ( .A(n960), .Y(n1007) );
  BUFX2 U67 ( .A(n960), .Y(n1006) );
  BUFX2 U68 ( .A(n959), .Y(n1004) );
  BUFX2 U69 ( .A(n959), .Y(n1003) );
  BUFX2 U70 ( .A(n958), .Y(n1001) );
  BUFX2 U71 ( .A(n958), .Y(n1000) );
  BUFX2 U72 ( .A(n957), .Y(n990) );
  BUFX2 U73 ( .A(n957), .Y(n989) );
  BUFX2 U74 ( .A(n956), .Y(n987) );
  BUFX2 U75 ( .A(n956), .Y(n986) );
  BUFX2 U76 ( .A(n955), .Y(n984) );
  BUFX2 U77 ( .A(n955), .Y(n983) );
  BUFX2 U78 ( .A(n954), .Y(n981) );
  BUFX2 U79 ( .A(n954), .Y(n980) );
  INVX1 U80 ( .A(\data_in_1c<0> ), .Y(n1028) );
  INVX1 U81 ( .A(\data_in_1c<1> ), .Y(n1029) );
  INVX1 U82 ( .A(\data_in_1c<2> ), .Y(n1030) );
  INVX1 U83 ( .A(\data_in_1c<3> ), .Y(n1031) );
  INVX1 U84 ( .A(\data_in_1c<4> ), .Y(n1032) );
  INVX1 U85 ( .A(\data_in_1c<5> ), .Y(n1033) );
  INVX1 U86 ( .A(\data_in_1c<6> ), .Y(n1034) );
  INVX1 U87 ( .A(\data_in_1c<7> ), .Y(n1035) );
  INVX1 U88 ( .A(\data_in_1c<8> ), .Y(n1036) );
  INVX1 U89 ( .A(\data_in_1c<9> ), .Y(n1037) );
  INVX1 U90 ( .A(\data_in_1c<10> ), .Y(n1038) );
  INVX1 U91 ( .A(\data_in_1c<11> ), .Y(n1039) );
  INVX1 U92 ( .A(\data_in_1c<12> ), .Y(n1040) );
  INVX1 U93 ( .A(\data_in_1c<13> ), .Y(n1041) );
  INVX1 U129 ( .A(\data_in_1c<14> ), .Y(n1042) );
  INVX1 U589 ( .A(\data_in_1c<15> ), .Y(n1043) );
  INVX1 U640 ( .A(wr), .Y(n1044) );
  INVX1 U659 ( .A(n1324), .Y(n1022) );
  INVX1 U660 ( .A(n1415), .Y(n1021) );
  INVX1 U664 ( .A(n1426), .Y(n1020) );
  INVX1 U666 ( .A(n1437), .Y(n1019) );
  INVX1 U672 ( .A(n1448), .Y(n1018) );
  INVX1 U675 ( .A(n1459), .Y(n1017) );
  INVX1 U679 ( .A(n1470), .Y(n1016) );
  INVX1 U682 ( .A(n1481), .Y(n1015) );
  AND2X1 U694 ( .A(wr1), .B(n1013), .Y(n1828) );
  INVX1 U697 ( .A(rst), .Y(n1013) );
  INVX2 U701 ( .A(n1013), .Y(n1012) );
  AND2X1 U706 ( .A(n387), .B(n372), .Y(n1) );
  INVX1 U712 ( .A(n1), .Y(n2) );
  AND2X1 U717 ( .A(n402), .B(n381), .Y(n3) );
  INVX1 U723 ( .A(n3), .Y(n4) );
  AND2X1 U728 ( .A(n1817), .B(n189), .Y(n5) );
  INVX1 U734 ( .A(n5), .Y(n6) );
  AND2X1 U739 ( .A(n973), .B(n289), .Y(n7) );
  INVX1 U745 ( .A(n7), .Y(n8) );
  OR2X1 U750 ( .A(n486), .B(n10), .Y(n9) );
  OR2X1 U756 ( .A(n473), .B(n474), .Y(n10) );
  OR2X1 U761 ( .A(n508), .B(n12), .Y(n11) );
  OR2X1 U767 ( .A(n487), .B(n507), .Y(n12) );
  OR2X1 U772 ( .A(n537), .B(n14), .Y(n13) );
  OR2X1 U786 ( .A(n522), .B(n523), .Y(n14) );
  OR2X1 U789 ( .A(n553), .B(n16), .Y(n15) );
  OR2X1 U801 ( .A(n538), .B(n552), .Y(n16) );
  OR2X1 U804 ( .A(n582), .B(n18), .Y(n17) );
  OR2X1 U816 ( .A(n567), .B(n568), .Y(n18) );
  OR2X1 U819 ( .A(n592), .B(n20), .Y(n19) );
  OR2X1 U831 ( .A(n583), .B(n591), .Y(n20) );
  OR2X1 U834 ( .A(n873), .B(n22), .Y(n21) );
  OR2X1 U846 ( .A(n871), .B(n872), .Y(n22) );
  OR2X1 U849 ( .A(n876), .B(n24), .Y(n23) );
  OR2X1 U861 ( .A(n874), .B(n875), .Y(n24) );
  OR2X1 U864 ( .A(n895), .B(n26), .Y(n25) );
  OR2X1 U870 ( .A(n893), .B(n894), .Y(n26) );
  OR2X1 U875 ( .A(n898), .B(n28), .Y(n27) );
  OR2X1 U882 ( .A(n896), .B(n897), .Y(n28) );
  OR2X1 U883 ( .A(n901), .B(n30), .Y(n29) );
  OR2X1 U884 ( .A(n899), .B(n900), .Y(n30) );
  OR2X1 U885 ( .A(n904), .B(n32), .Y(n31) );
  OR2X1 U886 ( .A(n902), .B(n903), .Y(n32) );
  OR2X1 U887 ( .A(n907), .B(n34), .Y(n33) );
  OR2X1 U888 ( .A(n905), .B(n906), .Y(n34) );
  OR2X1 U889 ( .A(n910), .B(n36), .Y(n35) );
  OR2X1 U890 ( .A(n908), .B(n909), .Y(n36) );
  OR2X1 U891 ( .A(n913), .B(n38), .Y(n37) );
  OR2X1 U892 ( .A(n911), .B(n912), .Y(n38) );
  OR2X1 U893 ( .A(n916), .B(n150), .Y(n50) );
  OR2X1 U894 ( .A(n914), .B(n915), .Y(n150) );
  AND2X1 U895 ( .A(n973), .B(n1828), .Y(n189) );
  AND2X1 U896 ( .A(n1828), .B(n1524), .Y(n289) );
  AND2X1 U897 ( .A(n940), .B(n942), .Y(n348) );
  INVX1 U898 ( .A(n348), .Y(n372) );
  AND2X1 U899 ( .A(n950), .B(n952), .Y(n379) );
  INVX1 U900 ( .A(n379), .Y(n381) );
  AND2X1 U901 ( .A(n940), .B(n941), .Y(n386) );
  INVX1 U902 ( .A(n386), .Y(n387) );
  AND2X1 U903 ( .A(n950), .B(n951), .Y(n401) );
  INVX1 U904 ( .A(n401), .Y(n402) );
  BUFX2 U905 ( .A(n1339), .Y(n408) );
  BUFX2 U906 ( .A(n1352), .Y(n409) );
  BUFX2 U907 ( .A(n1365), .Y(n421) );
  BUFX2 U908 ( .A(n1378), .Y(n422) );
  BUFX2 U909 ( .A(n1391), .Y(n434) );
  BUFX2 U910 ( .A(n1404), .Y(n435) );
  BUFX2 U911 ( .A(n1494), .Y(n447) );
  BUFX2 U912 ( .A(n1505), .Y(n448) );
  AND2X2 U913 ( .A(rd), .B(n1508), .Y(n460) );
  INVX1 U914 ( .A(n460), .Y(n461) );
  INVX1 U915 ( .A(n1314), .Y(n473) );
  INVX1 U916 ( .A(n1315), .Y(n474) );
  INVX1 U917 ( .A(n1316), .Y(n486) );
  INVX1 U918 ( .A(n1407), .Y(n487) );
  INVX1 U919 ( .A(n1408), .Y(n507) );
  INVX1 U920 ( .A(n1409), .Y(n508) );
  INVX1 U921 ( .A(n1418), .Y(n522) );
  INVX1 U922 ( .A(n1419), .Y(n523) );
  INVX1 U923 ( .A(n1420), .Y(n537) );
  INVX1 U924 ( .A(n1429), .Y(n538) );
  INVX1 U925 ( .A(n1430), .Y(n552) );
  INVX1 U926 ( .A(n1431), .Y(n553) );
  INVX1 U927 ( .A(n1440), .Y(n567) );
  INVX1 U928 ( .A(n1441), .Y(n568) );
  INVX1 U929 ( .A(n1442), .Y(n582) );
  INVX1 U930 ( .A(n1451), .Y(n583) );
  INVX1 U931 ( .A(n1452), .Y(n591) );
  INVX1 U932 ( .A(n1453), .Y(n592) );
  INVX1 U933 ( .A(n1462), .Y(n871) );
  INVX1 U934 ( .A(n1463), .Y(n872) );
  INVX1 U935 ( .A(n1464), .Y(n873) );
  INVX1 U936 ( .A(n1473), .Y(n874) );
  INVX1 U937 ( .A(n1474), .Y(n875) );
  INVX1 U938 ( .A(n1475), .Y(n876) );
  AND2X2 U939 ( .A(n1328), .B(n1327), .Y(n877) );
  INVX1 U940 ( .A(n877), .Y(n878) );
  AND2X2 U941 ( .A(n1341), .B(n1340), .Y(n879) );
  INVX1 U942 ( .A(n879), .Y(n880) );
  AND2X2 U943 ( .A(n1354), .B(n1353), .Y(n881) );
  INVX1 U944 ( .A(n881), .Y(n882) );
  AND2X2 U945 ( .A(n1367), .B(n1366), .Y(n883) );
  INVX1 U946 ( .A(n883), .Y(n884) );
  AND2X2 U947 ( .A(n1380), .B(n1379), .Y(n885) );
  INVX1 U948 ( .A(n885), .Y(n886) );
  AND2X2 U949 ( .A(n1393), .B(n1392), .Y(n887) );
  INVX1 U950 ( .A(n887), .Y(n888) );
  AND2X2 U951 ( .A(n1483), .B(n1482), .Y(n889) );
  INVX1 U952 ( .A(n889), .Y(n890) );
  AND2X2 U953 ( .A(n1496), .B(n1495), .Y(n891) );
  INVX1 U954 ( .A(n891), .Y(n892) );
  INVX1 U955 ( .A(n1321), .Y(n893) );
  INVX1 U956 ( .A(n1322), .Y(n894) );
  INVX1 U957 ( .A(n1323), .Y(n895) );
  INVX1 U958 ( .A(n1412), .Y(n896) );
  INVX1 U959 ( .A(n1413), .Y(n897) );
  INVX1 U960 ( .A(n1414), .Y(n898) );
  INVX1 U961 ( .A(n1423), .Y(n899) );
  INVX1 U962 ( .A(n1424), .Y(n900) );
  INVX1 U963 ( .A(n1425), .Y(n901) );
  INVX1 U964 ( .A(n1434), .Y(n902) );
  INVX1 U965 ( .A(n1435), .Y(n903) );
  INVX1 U966 ( .A(n1436), .Y(n904) );
  INVX1 U967 ( .A(n1445), .Y(n905) );
  INVX1 U968 ( .A(n1446), .Y(n906) );
  INVX1 U969 ( .A(n1447), .Y(n907) );
  INVX1 U970 ( .A(n1456), .Y(n908) );
  INVX1 U971 ( .A(n1457), .Y(n909) );
  INVX1 U972 ( .A(n1458), .Y(n910) );
  INVX1 U973 ( .A(n1467), .Y(n911) );
  INVX1 U974 ( .A(n1468), .Y(n912) );
  INVX1 U975 ( .A(n1469), .Y(n913) );
  INVX1 U976 ( .A(n1478), .Y(n914) );
  INVX1 U977 ( .A(n1479), .Y(n915) );
  INVX1 U978 ( .A(n1480), .Y(n916) );
  AND2X2 U979 ( .A(n1330), .B(n1329), .Y(n917) );
  INVX1 U980 ( .A(n917), .Y(n918) );
  AND2X2 U981 ( .A(n1343), .B(n1342), .Y(n919) );
  INVX1 U982 ( .A(n919), .Y(n920) );
  AND2X2 U983 ( .A(n1356), .B(n1355), .Y(n921) );
  INVX1 U984 ( .A(n921), .Y(n922) );
  AND2X2 U985 ( .A(n1369), .B(n1368), .Y(n923) );
  INVX1 U986 ( .A(n923), .Y(n924) );
  AND2X2 U987 ( .A(n1382), .B(n1381), .Y(n925) );
  INVX1 U988 ( .A(n925), .Y(n926) );
  AND2X2 U989 ( .A(n1395), .B(n1394), .Y(n927) );
  INVX1 U990 ( .A(n927), .Y(n928) );
  AND2X2 U991 ( .A(n1485), .B(n1484), .Y(n929) );
  INVX1 U992 ( .A(n929), .Y(n930) );
  AND2X2 U993 ( .A(n1498), .B(n1497), .Y(n931) );
  INVX1 U994 ( .A(n931), .Y(n932) );
  BUFX2 U995 ( .A(n1337), .Y(n933) );
  BUFX2 U996 ( .A(n1350), .Y(n934) );
  BUFX2 U997 ( .A(n1363), .Y(n935) );
  BUFX2 U998 ( .A(n1376), .Y(n936) );
  BUFX2 U999 ( .A(n1389), .Y(n937) );
  BUFX2 U1000 ( .A(n1402), .Y(n938) );
  BUFX2 U1001 ( .A(n1492), .Y(n939) );
  INVX1 U1002 ( .A(n970), .Y(n940) );
  INVX1 U1003 ( .A(n1499), .Y(n941) );
  INVX1 U1004 ( .A(n1500), .Y(n942) );
  BUFX2 U1005 ( .A(n1552), .Y(n970) );
  BUFX2 U1006 ( .A(n1335), .Y(n943) );
  BUFX2 U1007 ( .A(n1348), .Y(n944) );
  BUFX2 U1008 ( .A(n1361), .Y(n945) );
  BUFX2 U1009 ( .A(n1374), .Y(n946) );
  BUFX2 U1010 ( .A(n1387), .Y(n947) );
  BUFX2 U1011 ( .A(n1400), .Y(n948) );
  BUFX2 U1012 ( .A(n1490), .Y(n949) );
  INVX1 U1013 ( .A(n971), .Y(n950) );
  INVX1 U1014 ( .A(n1501), .Y(n951) );
  INVX1 U1015 ( .A(n1502), .Y(n952) );
  BUFX2 U1016 ( .A(n1514), .Y(n971) );
  BUFX2 U1017 ( .A(n1838), .Y(err) );
  BUFX2 U1018 ( .A(n1523), .Y(n972) );
  BUFX2 U1019 ( .A(n1541), .Y(n974) );
  BUFX2 U1020 ( .A(n1551), .Y(n975) );
  BUFX2 U1021 ( .A(n1561), .Y(n976) );
  BUFX2 U1022 ( .A(n1571), .Y(n977) );
  BUFX2 U1023 ( .A(n1580), .Y(n978) );
  BUFX2 U1024 ( .A(n1590), .Y(n979) );
  BUFX2 U1025 ( .A(n1610), .Y(n982) );
  BUFX2 U1026 ( .A(n1629), .Y(n985) );
  BUFX2 U1027 ( .A(n1650), .Y(n988) );
  BUFX2 U1028 ( .A(n1670), .Y(n991) );
  BUFX2 U1029 ( .A(n1679), .Y(n992) );
  BUFX2 U1030 ( .A(n1689), .Y(n993) );
  BUFX2 U1031 ( .A(n1698), .Y(n994) );
  BUFX2 U1032 ( .A(n1708), .Y(n995) );
  BUFX2 U1033 ( .A(n1717), .Y(n996) );
  BUFX2 U1034 ( .A(n1727), .Y(n997) );
  BUFX2 U1035 ( .A(n1736), .Y(n998) );
  BUFX2 U1036 ( .A(n1746), .Y(n999) );
  BUFX2 U1037 ( .A(n1765), .Y(n1002) );
  BUFX2 U1038 ( .A(n1785), .Y(n1005) );
  BUFX2 U1039 ( .A(n1805), .Y(n1008) );
  BUFX2 U1040 ( .A(n1818), .Y(n973) );
  AND2X1 U1041 ( .A(n1630), .B(n1318), .Y(n1817) );
  BUFX2 U1042 ( .A(n1837), .Y(n1011) );
  BUFX2 U1043 ( .A(n1600), .Y(n954) );
  BUFX2 U1044 ( .A(n1619), .Y(n955) );
  BUFX2 U1045 ( .A(n1640), .Y(n956) );
  BUFX2 U1046 ( .A(n1660), .Y(n957) );
  BUFX2 U1047 ( .A(n1755), .Y(n958) );
  BUFX2 U1048 ( .A(n1775), .Y(n959) );
  BUFX2 U1049 ( .A(n1795), .Y(n960) );
  BUFX2 U1050 ( .A(n1816), .Y(n961) );
  AND2X1 U1051 ( .A(enable), .B(n1013), .Y(n962) );
  INVX1 U1052 ( .A(n962), .Y(n963) );
  AND2X1 U1053 ( .A(n1513), .B(n1512), .Y(n964) );
  INVX1 U1054 ( .A(n964), .Y(n965) );
  INVX1 U1055 ( .A(n966), .Y(n967) );
  INVX1 U1056 ( .A(n968), .Y(n969) );
  AND2X1 U1057 ( .A(n950), .B(n1310), .Y(n1524) );
endmodule


module final_memory_0 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), err, .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<12> , \addr<11> , \addr<10> , \addr<9> , 
        \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , 
        \addr<2> , \addr<1> , \addr<0> }), wr, rd, enable, create_dump, 
    .bank_id({\bank_id<1> , \bank_id<0> }), clk, rst );
  input \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , \addr<12> , \addr<11> ,
         \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> , \addr<5> ,
         \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> , wr, rd, enable,
         create_dump, \bank_id<1> , \bank_id<0> , clk, rst;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , err;
  wire   n1838, rd0, wr0, rd1, wr1, \addr_1c<12> , \addr_1c<11> ,
         \addr_1c<10> , \addr_1c<9> , \addr_1c<8> , \addr_1c<7> , \addr_1c<6> ,
         \addr_1c<5> , \addr_1c<4> , \addr_1c<3> , \addr_1c<2> , \addr_1c<1> ,
         \addr_1c<0> , \data_in_1c<15> , \data_in_1c<14> , \data_in_1c<13> ,
         \data_in_1c<12> , \data_in_1c<11> , \data_in_1c<10> , \data_in_1c<9> ,
         \data_in_1c<8> , \data_in_1c<7> , \data_in_1c<6> , \data_in_1c<5> ,
         \data_in_1c<4> , \data_in_1c<3> , \data_in_1c<2> , \data_in_1c<1> ,
         \data_in_1c<0> , \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> ,
         \mem<0><3> , \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><7> ,
         \mem<1><6> , \mem<1><5> , \mem<1><4> , \mem<1><3> , \mem<1><2> ,
         \mem<1><1> , \mem<1><0> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><7> , \mem<3><6> , \mem<3><5> , \mem<3><4> , \mem<3><3> ,
         \mem<3><2> , \mem<3><1> , \mem<3><0> , \mem<4><7> , \mem<4><6> ,
         \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> , \mem<4><1> ,
         \mem<4><0> , \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> ,
         \mem<5><3> , \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><7> ,
         \mem<6><6> , \mem<6><5> , \mem<6><4> , \mem<6><3> , \mem<6><2> ,
         \mem<6><1> , \mem<6><0> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><7> , \mem<8><6> , \mem<8><5> , \mem<8><4> , \mem<8><3> ,
         \mem<8><2> , \mem<8><1> , \mem<8><0> , \mem<9><7> , \mem<9><6> ,
         \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> , \mem<9><1> ,
         \mem<9><0> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><7> ,
         \mem<11><6> , \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> ,
         \mem<11><1> , \mem<11><0> , \mem<12><7> , \mem<12><6> , \mem<12><5> ,
         \mem<12><4> , \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> ,
         \mem<13><7> , \mem<13><6> , \mem<13><5> , \mem<13><4> , \mem<13><3> ,
         \mem<13><2> , \mem<13><1> , \mem<13><0> , \mem<14><7> , \mem<14><6> ,
         \mem<14><5> , \mem<14><4> , \mem<14><3> , \mem<14><2> , \mem<14><1> ,
         \mem<14><0> , \mem<15><7> , \mem<15><6> , \mem<15><5> , \mem<15><4> ,
         \mem<15><3> , \mem<15><2> , \mem<15><1> , \mem<15><0> , \mem<16><7> ,
         \mem<16><6> , \mem<16><5> , \mem<16><4> , \mem<16><3> , \mem<16><2> ,
         \mem<16><1> , \mem<16><0> , \mem<17><7> , \mem<17><6> , \mem<17><5> ,
         \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> , \mem<17><0> ,
         \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> , \mem<18><3> ,
         \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><7> ,
         \mem<21><6> , \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> ,
         \mem<21><1> , \mem<21><0> , \mem<22><7> , \mem<22><6> , \mem<22><5> ,
         \mem<22><4> , \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> ,
         \mem<23><7> , \mem<23><6> , \mem<23><5> , \mem<23><4> , \mem<23><3> ,
         \mem<23><2> , \mem<23><1> , \mem<23><0> , \mem<24><7> , \mem<24><6> ,
         \mem<24><5> , \mem<24><4> , \mem<24><3> , \mem<24><2> , \mem<24><1> ,
         \mem<24><0> , \mem<25><7> , \mem<25><6> , \mem<25><5> , \mem<25><4> ,
         \mem<25><3> , \mem<25><2> , \mem<25><1> , \mem<25><0> , \mem<26><7> ,
         \mem<26><6> , \mem<26><5> , \mem<26><4> , \mem<26><3> , \mem<26><2> ,
         \mem<26><1> , \mem<26><0> , \mem<27><7> , \mem<27><6> , \mem<27><5> ,
         \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> , \mem<27><0> ,
         \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> , \mem<28><3> ,
         \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><7> ,
         \mem<31><6> , \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> ,
         \mem<31><1> , \mem<31><0> , \mem<32><7> , \mem<32><6> , \mem<32><5> ,
         \mem<32><4> , \mem<32><3> , \mem<32><2> , \mem<32><1> , \mem<32><0> ,
         \data_out_1c<15> , \data_out_1c<14> , \data_out_1c<13> ,
         \data_out_1c<12> , \data_out_1c<11> , \data_out_1c<10> ,
         \data_out_1c<9> , \data_out_1c<8> , rd2, wr2, rd3, wr3, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n50, n150, n189, n289, n348, n372, n379,
         n381, n386, n387, n401, n402, n408, n409, n421, n422, n434, n435,
         n447, n448, n460, n461, n473, n474, n486, n487, n507, n508, n522,
         n523, n537, n538, n552, n553, n567, n568, n582, n583, n591, n592,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837;

  DFFPOSX1 \mem_reg<0><7>  ( .D(n1046), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1047), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1048), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1049), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1050), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1051), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1052), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1053), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1054), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1055), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1056), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1057), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1058), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1059), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1060), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1061), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1062), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1063), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1064), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1065), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1066), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1067), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1068), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1069), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1070), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1071), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1072), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1073), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1074), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1075), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1076), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1077), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1078), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1079), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1080), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1081), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1082), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1083), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1084), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1085), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1086), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1087), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1088), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1089), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1090), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1091), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1092), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1093), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1094), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1095), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1096), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1097), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1098), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1099), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1100), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1101), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1102), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1103), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1104), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1105), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1106), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1107), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1108), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1109), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1110), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1111), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1112), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1113), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1114), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1115), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1116), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1117), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n1118), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n1119), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n1120), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n1121), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n1122), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n1123), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n1124), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n1125), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n1126), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n1127), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n1128), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n1129), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n1130), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n1131), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n1132), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n1133), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n1134), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n1135), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n1136), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n1137), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n1138), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n1139), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n1140), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n1141), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n1142), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n1143), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n1144), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n1145), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n1146), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n1147), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n1148), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n1149), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n1150), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n1151), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n1152), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n1153), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n1154), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n1155), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n1156), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n1157), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n1158), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n1159), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n1160), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n1161), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n1162), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n1163), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n1164), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n1165), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n1166), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n1167), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n1168), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n1169), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n1170), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n1171), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n1172), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n1173), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n1174), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n1175), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n1176), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n1177), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n1178), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n1179), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n1180), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n1181), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n1182), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n1183), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n1184), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n1185), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n1186), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n1187), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n1188), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n1189), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n1190), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n1191), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n1192), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n1193), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n1194), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n1195), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n1196), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n1197), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n1198), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n1199), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n1200), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n1201), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n1202), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n1203), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n1204), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n1205), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n1206), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n1207), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n1208), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n1209), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n1210), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n1211), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n1212), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n1213), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n1214), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n1215), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n1216), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n1217), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n1218), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n1219), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n1220), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n1221), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n1222), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n1223), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n1224), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n1225), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n1226), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n1227), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n1228), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n1229), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n1230), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n1231), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n1232), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n1233), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n1234), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n1235), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n1236), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n1237), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n1238), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n1239), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n1240), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n1241), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n1242), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n1243), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n1244), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n1245), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n1246), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n1247), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n1248), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n1249), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n1250), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n1251), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n1252), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n1253), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n1254), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n1255), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n1256), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n1257), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n1258), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n1259), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n1260), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n1261), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n1262), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n1263), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n1264), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n1265), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n1266), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n1267), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n1268), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n1269), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n1270), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n1271), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n1272), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n1273), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n1274), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n1275), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n1276), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n1277), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n1278), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n1279), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n1280), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n1281), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n1282), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n1283), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n1284), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n1285), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n1286), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n1287), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n1288), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n1289), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n1290), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n1291), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n1292), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n1293), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n1294), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n1295), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n1296), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n1297), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n1298), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n1299), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n1300), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n1301), .CLK(clk), .Q(\mem<31><0> ) );
  DFFPOSX1 \mem_reg<32><7>  ( .D(n1302), .CLK(clk), .Q(\mem<32><7> ) );
  DFFPOSX1 \mem_reg<32><6>  ( .D(n1303), .CLK(clk), .Q(\mem<32><6> ) );
  DFFPOSX1 \mem_reg<32><5>  ( .D(n1304), .CLK(clk), .Q(\mem<32><5> ) );
  DFFPOSX1 \mem_reg<32><4>  ( .D(n1305), .CLK(clk), .Q(\mem<32><4> ) );
  DFFPOSX1 \mem_reg<32><3>  ( .D(n1306), .CLK(clk), .Q(\mem<32><3> ) );
  DFFPOSX1 \mem_reg<32><2>  ( .D(n1307), .CLK(clk), .Q(\mem<32><2> ) );
  DFFPOSX1 \mem_reg<32><1>  ( .D(n1308), .CLK(clk), .Q(\mem<32><1> ) );
  DFFPOSX1 \mem_reg<32><0>  ( .D(n1309), .CLK(clk), .Q(\mem<32><0> ) );
  AND2X2 U9 ( .A(n1477), .B(n1476), .Y(n1478) );
  AND2X2 U10 ( .A(n1472), .B(n1471), .Y(n1473) );
  AND2X2 U11 ( .A(n1466), .B(n1465), .Y(n1467) );
  AND2X2 U12 ( .A(n1461), .B(n1460), .Y(n1462) );
  AND2X2 U13 ( .A(n1455), .B(n1454), .Y(n1456) );
  AND2X2 U14 ( .A(n1450), .B(n1449), .Y(n1451) );
  AND2X2 U15 ( .A(n1444), .B(n1443), .Y(n1445) );
  AND2X2 U16 ( .A(n1439), .B(n1438), .Y(n1440) );
  AND2X2 U17 ( .A(n1433), .B(n1432), .Y(n1434) );
  AND2X2 U18 ( .A(n1428), .B(n1427), .Y(n1429) );
  AND2X2 U19 ( .A(n1422), .B(n1421), .Y(n1423) );
  AND2X2 U20 ( .A(n1417), .B(n1416), .Y(n1418) );
  AND2X2 U21 ( .A(n1411), .B(n1410), .Y(n1412) );
  AND2X2 U22 ( .A(n1406), .B(n1405), .Y(n1407) );
  AND2X2 U30 ( .A(n1326), .B(n1024), .Y(n1631) );
  AND2X2 U31 ( .A(n1325), .B(n1024), .Y(n1786) );
  AND2X2 U32 ( .A(n1326), .B(\addr_1c<0> ), .Y(n1651) );
  AND2X2 U33 ( .A(n1325), .B(\addr_1c<0> ), .Y(n1806) );
  AND2X2 U34 ( .A(n1320), .B(n1319), .Y(n1321) );
  AND2X2 U45 ( .A(n1313), .B(n1312), .Y(n1314) );
  NOR3X1 U94 ( .A(n1044), .B(rd), .C(n963), .Y(wr0) );
  NOR3X1 U95 ( .A(n1045), .B(wr), .C(n963), .Y(rd0) );
  OAI21X1 U96 ( .A(n1011), .B(n1036), .C(n1836), .Y(n1309) );
  NAND2X1 U97 ( .A(\mem<32><0> ), .B(n1011), .Y(n1836) );
  OAI21X1 U98 ( .A(n1011), .B(n1037), .C(n1835), .Y(n1308) );
  NAND2X1 U99 ( .A(\mem<32><1> ), .B(n1011), .Y(n1835) );
  OAI21X1 U100 ( .A(n1011), .B(n1038), .C(n1834), .Y(n1307) );
  NAND2X1 U101 ( .A(\mem<32><2> ), .B(n1011), .Y(n1834) );
  OAI21X1 U102 ( .A(n1011), .B(n1039), .C(n1833), .Y(n1306) );
  NAND2X1 U103 ( .A(\mem<32><3> ), .B(n1011), .Y(n1833) );
  OAI21X1 U104 ( .A(n1011), .B(n1040), .C(n1832), .Y(n1305) );
  NAND2X1 U105 ( .A(\mem<32><4> ), .B(n1011), .Y(n1832) );
  OAI21X1 U106 ( .A(n1011), .B(n1041), .C(n1831), .Y(n1304) );
  NAND2X1 U107 ( .A(\mem<32><5> ), .B(n1011), .Y(n1831) );
  OAI21X1 U108 ( .A(n1011), .B(n1042), .C(n1830), .Y(n1303) );
  NAND2X1 U109 ( .A(\mem<32><6> ), .B(n1011), .Y(n1830) );
  OAI21X1 U110 ( .A(n1011), .B(n1043), .C(n1829), .Y(n1302) );
  NAND2X1 U111 ( .A(\mem<32><7> ), .B(n1011), .Y(n1829) );
  NAND3X1 U112 ( .A(n1828), .B(n1827), .C(n964), .Y(n1837) );
  OAI21X1 U113 ( .A(n6), .B(n1028), .C(n1826), .Y(n1301) );
  NAND2X1 U114 ( .A(\mem<31><0> ), .B(n6), .Y(n1826) );
  OAI21X1 U115 ( .A(n6), .B(n1029), .C(n1825), .Y(n1300) );
  NAND2X1 U116 ( .A(\mem<31><1> ), .B(n6), .Y(n1825) );
  OAI21X1 U117 ( .A(n6), .B(n1030), .C(n1824), .Y(n1299) );
  NAND2X1 U118 ( .A(\mem<31><2> ), .B(n6), .Y(n1824) );
  OAI21X1 U119 ( .A(n6), .B(n1031), .C(n1823), .Y(n1298) );
  NAND2X1 U120 ( .A(\mem<31><3> ), .B(n6), .Y(n1823) );
  OAI21X1 U121 ( .A(n6), .B(n1032), .C(n1822), .Y(n1297) );
  NAND2X1 U122 ( .A(\mem<31><4> ), .B(n6), .Y(n1822) );
  OAI21X1 U123 ( .A(n6), .B(n1033), .C(n1821), .Y(n1296) );
  NAND2X1 U124 ( .A(\mem<31><5> ), .B(n6), .Y(n1821) );
  OAI21X1 U125 ( .A(n6), .B(n1034), .C(n1820), .Y(n1295) );
  NAND2X1 U126 ( .A(\mem<31><6> ), .B(n6), .Y(n1820) );
  OAI21X1 U127 ( .A(n6), .B(n1035), .C(n1819), .Y(n1294) );
  NAND2X1 U128 ( .A(\mem<31><7> ), .B(n6), .Y(n1819) );
  OAI21X1 U130 ( .A(n1036), .B(n1010), .C(n1815), .Y(n1293) );
  NAND2X1 U131 ( .A(\mem<30><0> ), .B(n1010), .Y(n1815) );
  OAI21X1 U132 ( .A(n1037), .B(n1009), .C(n1814), .Y(n1292) );
  NAND2X1 U133 ( .A(\mem<30><1> ), .B(n1010), .Y(n1814) );
  OAI21X1 U134 ( .A(n1038), .B(n1009), .C(n1813), .Y(n1291) );
  NAND2X1 U135 ( .A(\mem<30><2> ), .B(n1010), .Y(n1813) );
  OAI21X1 U136 ( .A(n1039), .B(n1009), .C(n1812), .Y(n1290) );
  NAND2X1 U137 ( .A(\mem<30><3> ), .B(n1010), .Y(n1812) );
  OAI21X1 U138 ( .A(n1040), .B(n1009), .C(n1811), .Y(n1289) );
  NAND2X1 U139 ( .A(\mem<30><4> ), .B(n1010), .Y(n1811) );
  OAI21X1 U140 ( .A(n1041), .B(n1009), .C(n1810), .Y(n1288) );
  NAND2X1 U141 ( .A(\mem<30><5> ), .B(n1010), .Y(n1810) );
  OAI21X1 U142 ( .A(n1042), .B(n1009), .C(n1809), .Y(n1287) );
  NAND2X1 U143 ( .A(\mem<30><6> ), .B(n1010), .Y(n1809) );
  OAI21X1 U144 ( .A(n1043), .B(n1009), .C(n1808), .Y(n1286) );
  NAND2X1 U145 ( .A(\mem<30><7> ), .B(n1010), .Y(n1808) );
  NAND3X1 U146 ( .A(n1807), .B(n1828), .C(n1806), .Y(n1816) );
  OAI21X1 U147 ( .A(n1028), .B(n1008), .C(n1804), .Y(n1285) );
  NAND2X1 U148 ( .A(\mem<29><0> ), .B(n1008), .Y(n1804) );
  OAI21X1 U149 ( .A(n1029), .B(n1008), .C(n1803), .Y(n1284) );
  NAND2X1 U150 ( .A(\mem<29><1> ), .B(n1008), .Y(n1803) );
  OAI21X1 U151 ( .A(n1030), .B(n1008), .C(n1802), .Y(n1283) );
  NAND2X1 U152 ( .A(\mem<29><2> ), .B(n1008), .Y(n1802) );
  OAI21X1 U153 ( .A(n1031), .B(n1008), .C(n1801), .Y(n1282) );
  NAND2X1 U154 ( .A(\mem<29><3> ), .B(n1008), .Y(n1801) );
  OAI21X1 U155 ( .A(n1032), .B(n1008), .C(n1800), .Y(n1281) );
  NAND2X1 U156 ( .A(\mem<29><4> ), .B(n1008), .Y(n1800) );
  OAI21X1 U157 ( .A(n1033), .B(n1008), .C(n1799), .Y(n1280) );
  NAND2X1 U158 ( .A(\mem<29><5> ), .B(n1008), .Y(n1799) );
  OAI21X1 U159 ( .A(n1034), .B(n1008), .C(n1798), .Y(n1279) );
  NAND2X1 U160 ( .A(\mem<29><6> ), .B(n1008), .Y(n1798) );
  OAI21X1 U161 ( .A(n1035), .B(n1008), .C(n1797), .Y(n1278) );
  NAND2X1 U162 ( .A(\mem<29><7> ), .B(n1008), .Y(n1797) );
  NAND3X1 U163 ( .A(n973), .B(n1828), .C(n1796), .Y(n1805) );
  OAI21X1 U164 ( .A(n1036), .B(n1007), .C(n1794), .Y(n1277) );
  NAND2X1 U165 ( .A(\mem<28><0> ), .B(n1007), .Y(n1794) );
  OAI21X1 U166 ( .A(n1037), .B(n1006), .C(n1793), .Y(n1276) );
  NAND2X1 U167 ( .A(\mem<28><1> ), .B(n1007), .Y(n1793) );
  OAI21X1 U168 ( .A(n1038), .B(n1006), .C(n1792), .Y(n1275) );
  NAND2X1 U169 ( .A(\mem<28><2> ), .B(n1007), .Y(n1792) );
  OAI21X1 U170 ( .A(n1039), .B(n1006), .C(n1791), .Y(n1274) );
  NAND2X1 U171 ( .A(\mem<28><3> ), .B(n1007), .Y(n1791) );
  OAI21X1 U172 ( .A(n1040), .B(n1006), .C(n1790), .Y(n1273) );
  NAND2X1 U173 ( .A(\mem<28><4> ), .B(n1007), .Y(n1790) );
  OAI21X1 U174 ( .A(n1041), .B(n1006), .C(n1789), .Y(n1272) );
  NAND2X1 U175 ( .A(\mem<28><5> ), .B(n1007), .Y(n1789) );
  OAI21X1 U176 ( .A(n1042), .B(n1006), .C(n1788), .Y(n1271) );
  NAND2X1 U177 ( .A(\mem<28><6> ), .B(n1007), .Y(n1788) );
  OAI21X1 U178 ( .A(n1043), .B(n1006), .C(n1787), .Y(n1270) );
  NAND2X1 U179 ( .A(\mem<28><7> ), .B(n1007), .Y(n1787) );
  NAND3X1 U180 ( .A(n1807), .B(n1828), .C(n1786), .Y(n1795) );
  OAI21X1 U181 ( .A(n1028), .B(n1005), .C(n1784), .Y(n1269) );
  NAND2X1 U182 ( .A(\mem<27><0> ), .B(n1005), .Y(n1784) );
  OAI21X1 U183 ( .A(n1029), .B(n1005), .C(n1783), .Y(n1268) );
  NAND2X1 U184 ( .A(\mem<27><1> ), .B(n1005), .Y(n1783) );
  OAI21X1 U185 ( .A(n1030), .B(n1005), .C(n1782), .Y(n1267) );
  NAND2X1 U186 ( .A(\mem<27><2> ), .B(n1005), .Y(n1782) );
  OAI21X1 U187 ( .A(n1031), .B(n1005), .C(n1781), .Y(n1266) );
  NAND2X1 U188 ( .A(\mem<27><3> ), .B(n1005), .Y(n1781) );
  OAI21X1 U189 ( .A(n1032), .B(n1005), .C(n1780), .Y(n1265) );
  NAND2X1 U190 ( .A(\mem<27><4> ), .B(n1005), .Y(n1780) );
  OAI21X1 U191 ( .A(n1033), .B(n1005), .C(n1779), .Y(n1264) );
  NAND2X1 U192 ( .A(\mem<27><5> ), .B(n1005), .Y(n1779) );
  OAI21X1 U193 ( .A(n1034), .B(n1005), .C(n1778), .Y(n1263) );
  NAND2X1 U194 ( .A(\mem<27><6> ), .B(n1005), .Y(n1778) );
  OAI21X1 U195 ( .A(n1035), .B(n1005), .C(n1777), .Y(n1262) );
  NAND2X1 U196 ( .A(\mem<27><7> ), .B(n1005), .Y(n1777) );
  NAND3X1 U197 ( .A(n973), .B(n1828), .C(n1776), .Y(n1785) );
  OAI21X1 U198 ( .A(n1036), .B(n1004), .C(n1774), .Y(n1261) );
  NAND2X1 U199 ( .A(\mem<26><0> ), .B(n1004), .Y(n1774) );
  OAI21X1 U200 ( .A(n1037), .B(n1003), .C(n1773), .Y(n1260) );
  NAND2X1 U201 ( .A(\mem<26><1> ), .B(n1004), .Y(n1773) );
  OAI21X1 U202 ( .A(n1038), .B(n1003), .C(n1772), .Y(n1259) );
  NAND2X1 U203 ( .A(\mem<26><2> ), .B(n1004), .Y(n1772) );
  OAI21X1 U204 ( .A(n1039), .B(n1003), .C(n1771), .Y(n1258) );
  NAND2X1 U205 ( .A(\mem<26><3> ), .B(n1004), .Y(n1771) );
  OAI21X1 U206 ( .A(n1040), .B(n1003), .C(n1770), .Y(n1257) );
  NAND2X1 U207 ( .A(\mem<26><4> ), .B(n1004), .Y(n1770) );
  OAI21X1 U208 ( .A(n1041), .B(n1003), .C(n1769), .Y(n1256) );
  NAND2X1 U209 ( .A(\mem<26><5> ), .B(n1004), .Y(n1769) );
  OAI21X1 U210 ( .A(n1042), .B(n1003), .C(n1768), .Y(n1255) );
  NAND2X1 U211 ( .A(\mem<26><6> ), .B(n1004), .Y(n1768) );
  OAI21X1 U212 ( .A(n1043), .B(n1003), .C(n1767), .Y(n1254) );
  NAND2X1 U213 ( .A(\mem<26><7> ), .B(n1004), .Y(n1767) );
  NAND3X1 U214 ( .A(n1806), .B(n1828), .C(n1766), .Y(n1775) );
  OAI21X1 U215 ( .A(n1028), .B(n1002), .C(n1764), .Y(n1253) );
  NAND2X1 U216 ( .A(\mem<25><0> ), .B(n1002), .Y(n1764) );
  OAI21X1 U217 ( .A(n1029), .B(n1002), .C(n1763), .Y(n1252) );
  NAND2X1 U218 ( .A(\mem<25><1> ), .B(n1002), .Y(n1763) );
  OAI21X1 U219 ( .A(n1030), .B(n1002), .C(n1762), .Y(n1251) );
  NAND2X1 U220 ( .A(\mem<25><2> ), .B(n1002), .Y(n1762) );
  OAI21X1 U221 ( .A(n1031), .B(n1002), .C(n1761), .Y(n1250) );
  NAND2X1 U222 ( .A(\mem<25><3> ), .B(n1002), .Y(n1761) );
  OAI21X1 U223 ( .A(n1032), .B(n1002), .C(n1760), .Y(n1249) );
  NAND2X1 U224 ( .A(\mem<25><4> ), .B(n1002), .Y(n1760) );
  OAI21X1 U225 ( .A(n1033), .B(n1002), .C(n1759), .Y(n1248) );
  NAND2X1 U226 ( .A(\mem<25><5> ), .B(n1002), .Y(n1759) );
  OAI21X1 U227 ( .A(n1034), .B(n1002), .C(n1758), .Y(n1247) );
  NAND2X1 U228 ( .A(\mem<25><6> ), .B(n1002), .Y(n1758) );
  OAI21X1 U229 ( .A(n1035), .B(n1002), .C(n1757), .Y(n1246) );
  NAND2X1 U230 ( .A(\mem<25><7> ), .B(n1002), .Y(n1757) );
  NAND3X1 U231 ( .A(n973), .B(n1828), .C(n1756), .Y(n1765) );
  OAI21X1 U232 ( .A(n1036), .B(n1001), .C(n1754), .Y(n1245) );
  NAND2X1 U233 ( .A(\mem<24><0> ), .B(n1001), .Y(n1754) );
  OAI21X1 U234 ( .A(n1037), .B(n1000), .C(n1753), .Y(n1244) );
  NAND2X1 U235 ( .A(\mem<24><1> ), .B(n1001), .Y(n1753) );
  OAI21X1 U236 ( .A(n1038), .B(n1000), .C(n1752), .Y(n1243) );
  NAND2X1 U237 ( .A(\mem<24><2> ), .B(n1001), .Y(n1752) );
  OAI21X1 U238 ( .A(n1039), .B(n1000), .C(n1751), .Y(n1242) );
  NAND2X1 U239 ( .A(\mem<24><3> ), .B(n1001), .Y(n1751) );
  OAI21X1 U240 ( .A(n1040), .B(n1000), .C(n1750), .Y(n1241) );
  NAND2X1 U241 ( .A(\mem<24><4> ), .B(n1001), .Y(n1750) );
  OAI21X1 U242 ( .A(n1041), .B(n1000), .C(n1749), .Y(n1240) );
  NAND2X1 U243 ( .A(\mem<24><5> ), .B(n1001), .Y(n1749) );
  OAI21X1 U244 ( .A(n1042), .B(n1000), .C(n1748), .Y(n1239) );
  NAND2X1 U245 ( .A(\mem<24><6> ), .B(n1001), .Y(n1748) );
  OAI21X1 U246 ( .A(n1043), .B(n1000), .C(n1747), .Y(n1238) );
  NAND2X1 U247 ( .A(\mem<24><7> ), .B(n1001), .Y(n1747) );
  NAND3X1 U248 ( .A(n1786), .B(n1828), .C(n1766), .Y(n1755) );
  OAI21X1 U249 ( .A(n1028), .B(n999), .C(n1745), .Y(n1237) );
  NAND2X1 U250 ( .A(\mem<23><0> ), .B(n999), .Y(n1745) );
  OAI21X1 U251 ( .A(n1029), .B(n999), .C(n1744), .Y(n1236) );
  NAND2X1 U252 ( .A(\mem<23><1> ), .B(n999), .Y(n1744) );
  OAI21X1 U253 ( .A(n1030), .B(n999), .C(n1743), .Y(n1235) );
  NAND2X1 U254 ( .A(\mem<23><2> ), .B(n999), .Y(n1743) );
  OAI21X1 U255 ( .A(n1031), .B(n999), .C(n1742), .Y(n1234) );
  NAND2X1 U256 ( .A(\mem<23><3> ), .B(n999), .Y(n1742) );
  OAI21X1 U257 ( .A(n1032), .B(n999), .C(n1741), .Y(n1233) );
  NAND2X1 U258 ( .A(\mem<23><4> ), .B(n999), .Y(n1741) );
  OAI21X1 U259 ( .A(n1033), .B(n999), .C(n1740), .Y(n1232) );
  NAND2X1 U260 ( .A(\mem<23><5> ), .B(n999), .Y(n1740) );
  OAI21X1 U261 ( .A(n1034), .B(n999), .C(n1739), .Y(n1231) );
  NAND2X1 U262 ( .A(\mem<23><6> ), .B(n999), .Y(n1739) );
  OAI21X1 U263 ( .A(n1035), .B(n999), .C(n1738), .Y(n1230) );
  NAND2X1 U264 ( .A(\mem<23><7> ), .B(n999), .Y(n1738) );
  NAND3X1 U265 ( .A(n973), .B(n1828), .C(n1737), .Y(n1746) );
  OAI21X1 U266 ( .A(n1036), .B(n998), .C(n1735), .Y(n1229) );
  NAND2X1 U267 ( .A(\mem<22><0> ), .B(n998), .Y(n1735) );
  OAI21X1 U268 ( .A(n1037), .B(n998), .C(n1734), .Y(n1228) );
  NAND2X1 U269 ( .A(\mem<22><1> ), .B(n998), .Y(n1734) );
  OAI21X1 U270 ( .A(n1038), .B(n998), .C(n1733), .Y(n1227) );
  NAND2X1 U271 ( .A(\mem<22><2> ), .B(n998), .Y(n1733) );
  OAI21X1 U272 ( .A(n1039), .B(n998), .C(n1732), .Y(n1226) );
  NAND2X1 U273 ( .A(\mem<22><3> ), .B(n998), .Y(n1732) );
  OAI21X1 U274 ( .A(n1040), .B(n998), .C(n1731), .Y(n1225) );
  NAND2X1 U275 ( .A(\mem<22><4> ), .B(n998), .Y(n1731) );
  OAI21X1 U276 ( .A(n1041), .B(n998), .C(n1730), .Y(n1224) );
  NAND2X1 U277 ( .A(\mem<22><5> ), .B(n998), .Y(n1730) );
  OAI21X1 U278 ( .A(n1042), .B(n998), .C(n1729), .Y(n1223) );
  NAND2X1 U279 ( .A(\mem<22><6> ), .B(n998), .Y(n1729) );
  OAI21X1 U280 ( .A(n1043), .B(n998), .C(n1728), .Y(n1222) );
  NAND2X1 U281 ( .A(\mem<22><7> ), .B(n998), .Y(n1728) );
  NAND3X1 U282 ( .A(n1806), .B(n1828), .C(n969), .Y(n1736) );
  OAI21X1 U283 ( .A(n1028), .B(n997), .C(n1726), .Y(n1221) );
  NAND2X1 U284 ( .A(\mem<21><0> ), .B(n997), .Y(n1726) );
  OAI21X1 U285 ( .A(n1029), .B(n997), .C(n1725), .Y(n1220) );
  NAND2X1 U286 ( .A(\mem<21><1> ), .B(n997), .Y(n1725) );
  OAI21X1 U287 ( .A(n1030), .B(n997), .C(n1724), .Y(n1219) );
  NAND2X1 U288 ( .A(\mem<21><2> ), .B(n997), .Y(n1724) );
  OAI21X1 U289 ( .A(n1031), .B(n997), .C(n1723), .Y(n1218) );
  NAND2X1 U290 ( .A(\mem<21><3> ), .B(n997), .Y(n1723) );
  OAI21X1 U291 ( .A(n1032), .B(n997), .C(n1722), .Y(n1217) );
  NAND2X1 U292 ( .A(\mem<21><4> ), .B(n997), .Y(n1722) );
  OAI21X1 U293 ( .A(n1033), .B(n997), .C(n1721), .Y(n1216) );
  NAND2X1 U294 ( .A(\mem<21><5> ), .B(n997), .Y(n1721) );
  OAI21X1 U295 ( .A(n1034), .B(n997), .C(n1720), .Y(n1215) );
  NAND2X1 U296 ( .A(\mem<21><6> ), .B(n997), .Y(n1720) );
  OAI21X1 U297 ( .A(n1035), .B(n997), .C(n1719), .Y(n1214) );
  NAND2X1 U298 ( .A(\mem<21><7> ), .B(n997), .Y(n1719) );
  NAND3X1 U299 ( .A(n973), .B(n1828), .C(n1718), .Y(n1727) );
  OAI21X1 U300 ( .A(n1036), .B(n996), .C(n1716), .Y(n1213) );
  NAND2X1 U301 ( .A(\mem<20><0> ), .B(n996), .Y(n1716) );
  OAI21X1 U302 ( .A(n1037), .B(n996), .C(n1715), .Y(n1212) );
  NAND2X1 U303 ( .A(\mem<20><1> ), .B(n996), .Y(n1715) );
  OAI21X1 U304 ( .A(n1038), .B(n996), .C(n1714), .Y(n1211) );
  NAND2X1 U305 ( .A(\mem<20><2> ), .B(n996), .Y(n1714) );
  OAI21X1 U306 ( .A(n1039), .B(n996), .C(n1713), .Y(n1210) );
  NAND2X1 U307 ( .A(\mem<20><3> ), .B(n996), .Y(n1713) );
  OAI21X1 U308 ( .A(n1040), .B(n996), .C(n1712), .Y(n1209) );
  NAND2X1 U309 ( .A(\mem<20><4> ), .B(n996), .Y(n1712) );
  OAI21X1 U310 ( .A(n1041), .B(n996), .C(n1711), .Y(n1208) );
  NAND2X1 U311 ( .A(\mem<20><5> ), .B(n996), .Y(n1711) );
  OAI21X1 U312 ( .A(n1042), .B(n996), .C(n1710), .Y(n1207) );
  NAND2X1 U313 ( .A(\mem<20><6> ), .B(n996), .Y(n1710) );
  OAI21X1 U314 ( .A(n1043), .B(n996), .C(n1709), .Y(n1206) );
  NAND2X1 U315 ( .A(\mem<20><7> ), .B(n996), .Y(n1709) );
  NAND3X1 U316 ( .A(n1786), .B(n1828), .C(n969), .Y(n1717) );
  OAI21X1 U317 ( .A(n1028), .B(n995), .C(n1707), .Y(n1205) );
  NAND2X1 U318 ( .A(\mem<19><0> ), .B(n995), .Y(n1707) );
  OAI21X1 U319 ( .A(n1029), .B(n995), .C(n1706), .Y(n1204) );
  NAND2X1 U320 ( .A(\mem<19><1> ), .B(n995), .Y(n1706) );
  OAI21X1 U321 ( .A(n1030), .B(n995), .C(n1705), .Y(n1203) );
  NAND2X1 U322 ( .A(\mem<19><2> ), .B(n995), .Y(n1705) );
  OAI21X1 U323 ( .A(n1031), .B(n995), .C(n1704), .Y(n1202) );
  NAND2X1 U324 ( .A(\mem<19><3> ), .B(n995), .Y(n1704) );
  OAI21X1 U325 ( .A(n1032), .B(n995), .C(n1703), .Y(n1201) );
  NAND2X1 U326 ( .A(\mem<19><4> ), .B(n995), .Y(n1703) );
  OAI21X1 U327 ( .A(n1033), .B(n995), .C(n1702), .Y(n1200) );
  NAND2X1 U328 ( .A(\mem<19><5> ), .B(n995), .Y(n1702) );
  OAI21X1 U329 ( .A(n1034), .B(n995), .C(n1701), .Y(n1199) );
  NAND2X1 U330 ( .A(\mem<19><6> ), .B(n995), .Y(n1701) );
  OAI21X1 U331 ( .A(n1035), .B(n995), .C(n1700), .Y(n1198) );
  NAND2X1 U332 ( .A(\mem<19><7> ), .B(n995), .Y(n1700) );
  NAND3X1 U333 ( .A(n973), .B(n1828), .C(n1699), .Y(n1708) );
  OAI21X1 U334 ( .A(n1036), .B(n994), .C(n1697), .Y(n1197) );
  NAND2X1 U335 ( .A(\mem<18><0> ), .B(n994), .Y(n1697) );
  OAI21X1 U336 ( .A(n1037), .B(n994), .C(n1696), .Y(n1196) );
  NAND2X1 U337 ( .A(\mem<18><1> ), .B(n994), .Y(n1696) );
  OAI21X1 U338 ( .A(n1038), .B(n994), .C(n1695), .Y(n1195) );
  NAND2X1 U339 ( .A(\mem<18><2> ), .B(n994), .Y(n1695) );
  OAI21X1 U340 ( .A(n1039), .B(n994), .C(n1694), .Y(n1194) );
  NAND2X1 U341 ( .A(\mem<18><3> ), .B(n994), .Y(n1694) );
  OAI21X1 U342 ( .A(n1040), .B(n994), .C(n1693), .Y(n1193) );
  NAND2X1 U343 ( .A(\mem<18><4> ), .B(n994), .Y(n1693) );
  OAI21X1 U344 ( .A(n1041), .B(n994), .C(n1692), .Y(n1192) );
  NAND2X1 U345 ( .A(\mem<18><5> ), .B(n994), .Y(n1692) );
  OAI21X1 U346 ( .A(n1042), .B(n994), .C(n1691), .Y(n1191) );
  NAND2X1 U347 ( .A(\mem<18><6> ), .B(n994), .Y(n1691) );
  OAI21X1 U348 ( .A(n1043), .B(n994), .C(n1690), .Y(n1190) );
  NAND2X1 U349 ( .A(\mem<18><7> ), .B(n994), .Y(n1690) );
  NAND3X1 U350 ( .A(n1806), .B(n1828), .C(n967), .Y(n1698) );
  OAI21X1 U351 ( .A(n1028), .B(n993), .C(n1688), .Y(n1189) );
  NAND2X1 U352 ( .A(\mem<17><0> ), .B(n993), .Y(n1688) );
  OAI21X1 U353 ( .A(n1029), .B(n993), .C(n1687), .Y(n1188) );
  NAND2X1 U354 ( .A(\mem<17><1> ), .B(n993), .Y(n1687) );
  OAI21X1 U355 ( .A(n1030), .B(n993), .C(n1686), .Y(n1187) );
  NAND2X1 U356 ( .A(\mem<17><2> ), .B(n993), .Y(n1686) );
  OAI21X1 U357 ( .A(n1031), .B(n993), .C(n1685), .Y(n1186) );
  NAND2X1 U358 ( .A(\mem<17><3> ), .B(n993), .Y(n1685) );
  OAI21X1 U359 ( .A(n1032), .B(n993), .C(n1684), .Y(n1185) );
  NAND2X1 U360 ( .A(\mem<17><4> ), .B(n993), .Y(n1684) );
  OAI21X1 U361 ( .A(n1033), .B(n993), .C(n1683), .Y(n1184) );
  NAND2X1 U362 ( .A(\mem<17><5> ), .B(n993), .Y(n1683) );
  OAI21X1 U363 ( .A(n1034), .B(n993), .C(n1682), .Y(n1183) );
  NAND2X1 U364 ( .A(\mem<17><6> ), .B(n993), .Y(n1682) );
  OAI21X1 U365 ( .A(n1035), .B(n993), .C(n1681), .Y(n1182) );
  NAND2X1 U366 ( .A(\mem<17><7> ), .B(n993), .Y(n1681) );
  NAND3X1 U367 ( .A(n973), .B(n1828), .C(n1680), .Y(n1689) );
  OAI21X1 U368 ( .A(n1036), .B(n992), .C(n1678), .Y(n1181) );
  NAND2X1 U369 ( .A(\mem<16><0> ), .B(n992), .Y(n1678) );
  OAI21X1 U370 ( .A(n1037), .B(n992), .C(n1677), .Y(n1180) );
  NAND2X1 U371 ( .A(\mem<16><1> ), .B(n992), .Y(n1677) );
  OAI21X1 U372 ( .A(n1038), .B(n992), .C(n1676), .Y(n1179) );
  NAND2X1 U373 ( .A(\mem<16><2> ), .B(n992), .Y(n1676) );
  OAI21X1 U374 ( .A(n1039), .B(n992), .C(n1675), .Y(n1178) );
  NAND2X1 U375 ( .A(\mem<16><3> ), .B(n992), .Y(n1675) );
  OAI21X1 U376 ( .A(n1040), .B(n992), .C(n1674), .Y(n1177) );
  NAND2X1 U377 ( .A(\mem<16><4> ), .B(n992), .Y(n1674) );
  OAI21X1 U378 ( .A(n1041), .B(n992), .C(n1673), .Y(n1176) );
  NAND2X1 U379 ( .A(\mem<16><5> ), .B(n992), .Y(n1673) );
  OAI21X1 U380 ( .A(n1042), .B(n992), .C(n1672), .Y(n1175) );
  NAND2X1 U381 ( .A(\mem<16><6> ), .B(n992), .Y(n1672) );
  OAI21X1 U382 ( .A(n1043), .B(n992), .C(n1671), .Y(n1174) );
  NAND2X1 U383 ( .A(\mem<16><7> ), .B(n992), .Y(n1671) );
  NAND3X1 U384 ( .A(n1786), .B(n1828), .C(n967), .Y(n1679) );
  OAI21X1 U385 ( .A(n1028), .B(n991), .C(n1669), .Y(n1173) );
  NAND2X1 U386 ( .A(\mem<15><0> ), .B(n991), .Y(n1669) );
  OAI21X1 U387 ( .A(n1029), .B(n991), .C(n1668), .Y(n1172) );
  NAND2X1 U388 ( .A(\mem<15><1> ), .B(n991), .Y(n1668) );
  OAI21X1 U389 ( .A(n1030), .B(n991), .C(n1667), .Y(n1171) );
  NAND2X1 U390 ( .A(\mem<15><2> ), .B(n991), .Y(n1667) );
  OAI21X1 U391 ( .A(n1031), .B(n991), .C(n1666), .Y(n1170) );
  NAND2X1 U392 ( .A(\mem<15><3> ), .B(n991), .Y(n1666) );
  OAI21X1 U393 ( .A(n1032), .B(n991), .C(n1665), .Y(n1169) );
  NAND2X1 U394 ( .A(\mem<15><4> ), .B(n991), .Y(n1665) );
  OAI21X1 U395 ( .A(n1033), .B(n991), .C(n1664), .Y(n1168) );
  NAND2X1 U396 ( .A(\mem<15><5> ), .B(n991), .Y(n1664) );
  OAI21X1 U397 ( .A(n1034), .B(n991), .C(n1663), .Y(n1167) );
  NAND2X1 U398 ( .A(\mem<15><6> ), .B(n991), .Y(n1663) );
  OAI21X1 U399 ( .A(n1035), .B(n991), .C(n1662), .Y(n1166) );
  NAND2X1 U400 ( .A(\mem<15><7> ), .B(n991), .Y(n1662) );
  NAND3X1 U401 ( .A(n973), .B(n1828), .C(n1661), .Y(n1670) );
  OAI21X1 U402 ( .A(n1036), .B(n990), .C(n1659), .Y(n1165) );
  NAND2X1 U403 ( .A(\mem<14><0> ), .B(n990), .Y(n1659) );
  OAI21X1 U404 ( .A(n1037), .B(n989), .C(n1658), .Y(n1164) );
  NAND2X1 U405 ( .A(\mem<14><1> ), .B(n990), .Y(n1658) );
  OAI21X1 U406 ( .A(n1038), .B(n989), .C(n1657), .Y(n1163) );
  NAND2X1 U407 ( .A(\mem<14><2> ), .B(n990), .Y(n1657) );
  OAI21X1 U408 ( .A(n1039), .B(n989), .C(n1656), .Y(n1162) );
  NAND2X1 U409 ( .A(\mem<14><3> ), .B(n990), .Y(n1656) );
  OAI21X1 U410 ( .A(n1040), .B(n989), .C(n1655), .Y(n1161) );
  NAND2X1 U411 ( .A(\mem<14><4> ), .B(n990), .Y(n1655) );
  OAI21X1 U412 ( .A(n1041), .B(n989), .C(n1654), .Y(n1160) );
  NAND2X1 U413 ( .A(\mem<14><5> ), .B(n990), .Y(n1654) );
  OAI21X1 U414 ( .A(n1042), .B(n989), .C(n1653), .Y(n1159) );
  NAND2X1 U415 ( .A(\mem<14><6> ), .B(n990), .Y(n1653) );
  OAI21X1 U416 ( .A(n1043), .B(n989), .C(n1652), .Y(n1158) );
  NAND2X1 U417 ( .A(\mem<14><7> ), .B(n990), .Y(n1652) );
  NAND3X1 U418 ( .A(n1807), .B(n1828), .C(n1651), .Y(n1660) );
  OAI21X1 U419 ( .A(n1028), .B(n988), .C(n1649), .Y(n1157) );
  NAND2X1 U420 ( .A(\mem<13><0> ), .B(n988), .Y(n1649) );
  OAI21X1 U421 ( .A(n1029), .B(n988), .C(n1648), .Y(n1156) );
  NAND2X1 U422 ( .A(\mem<13><1> ), .B(n988), .Y(n1648) );
  OAI21X1 U423 ( .A(n1030), .B(n988), .C(n1647), .Y(n1155) );
  NAND2X1 U424 ( .A(\mem<13><2> ), .B(n988), .Y(n1647) );
  OAI21X1 U425 ( .A(n1031), .B(n988), .C(n1646), .Y(n1154) );
  NAND2X1 U426 ( .A(\mem<13><3> ), .B(n988), .Y(n1646) );
  OAI21X1 U427 ( .A(n1032), .B(n988), .C(n1645), .Y(n1153) );
  NAND2X1 U428 ( .A(\mem<13><4> ), .B(n988), .Y(n1645) );
  OAI21X1 U429 ( .A(n1033), .B(n988), .C(n1644), .Y(n1152) );
  NAND2X1 U430 ( .A(\mem<13><5> ), .B(n988), .Y(n1644) );
  OAI21X1 U431 ( .A(n1034), .B(n988), .C(n1643), .Y(n1151) );
  NAND2X1 U432 ( .A(\mem<13><6> ), .B(n988), .Y(n1643) );
  OAI21X1 U433 ( .A(n1035), .B(n988), .C(n1642), .Y(n1150) );
  NAND2X1 U434 ( .A(\mem<13><7> ), .B(n988), .Y(n1642) );
  NAND3X1 U435 ( .A(n973), .B(n1828), .C(n1641), .Y(n1650) );
  OAI21X1 U436 ( .A(n1036), .B(n987), .C(n1639), .Y(n1149) );
  NAND2X1 U437 ( .A(\mem<12><0> ), .B(n987), .Y(n1639) );
  OAI21X1 U438 ( .A(n1037), .B(n986), .C(n1638), .Y(n1148) );
  NAND2X1 U439 ( .A(\mem<12><1> ), .B(n987), .Y(n1638) );
  OAI21X1 U440 ( .A(n1038), .B(n986), .C(n1637), .Y(n1147) );
  NAND2X1 U441 ( .A(\mem<12><2> ), .B(n987), .Y(n1637) );
  OAI21X1 U442 ( .A(n1039), .B(n986), .C(n1636), .Y(n1146) );
  NAND2X1 U443 ( .A(\mem<12><3> ), .B(n987), .Y(n1636) );
  OAI21X1 U444 ( .A(n1040), .B(n986), .C(n1635), .Y(n1145) );
  NAND2X1 U445 ( .A(\mem<12><4> ), .B(n987), .Y(n1635) );
  OAI21X1 U446 ( .A(n1041), .B(n986), .C(n1634), .Y(n1144) );
  NAND2X1 U447 ( .A(\mem<12><5> ), .B(n987), .Y(n1634) );
  OAI21X1 U448 ( .A(n1042), .B(n986), .C(n1633), .Y(n1143) );
  NAND2X1 U449 ( .A(\mem<12><6> ), .B(n987), .Y(n1633) );
  OAI21X1 U450 ( .A(n1043), .B(n986), .C(n1632), .Y(n1142) );
  NAND2X1 U451 ( .A(\mem<12><7> ), .B(n987), .Y(n1632) );
  NAND3X1 U452 ( .A(n1807), .B(n1828), .C(n1631), .Y(n1640) );
  OAI21X1 U453 ( .A(n1028), .B(n985), .C(n1628), .Y(n1141) );
  NAND2X1 U454 ( .A(\mem<11><0> ), .B(n985), .Y(n1628) );
  OAI21X1 U455 ( .A(n1029), .B(n985), .C(n1627), .Y(n1140) );
  NAND2X1 U456 ( .A(\mem<11><1> ), .B(n985), .Y(n1627) );
  OAI21X1 U457 ( .A(n1030), .B(n985), .C(n1626), .Y(n1139) );
  NAND2X1 U458 ( .A(\mem<11><2> ), .B(n985), .Y(n1626) );
  OAI21X1 U459 ( .A(n1031), .B(n985), .C(n1625), .Y(n1138) );
  NAND2X1 U460 ( .A(\mem<11><3> ), .B(n985), .Y(n1625) );
  OAI21X1 U461 ( .A(n1032), .B(n985), .C(n1624), .Y(n1137) );
  NAND2X1 U462 ( .A(\mem<11><4> ), .B(n985), .Y(n1624) );
  OAI21X1 U463 ( .A(n1033), .B(n985), .C(n1623), .Y(n1136) );
  NAND2X1 U464 ( .A(\mem<11><5> ), .B(n985), .Y(n1623) );
  OAI21X1 U465 ( .A(n1034), .B(n985), .C(n1622), .Y(n1135) );
  NAND2X1 U466 ( .A(\mem<11><6> ), .B(n985), .Y(n1622) );
  OAI21X1 U467 ( .A(n1035), .B(n985), .C(n1621), .Y(n1134) );
  NAND2X1 U468 ( .A(\mem<11><7> ), .B(n985), .Y(n1621) );
  NAND3X1 U469 ( .A(n973), .B(n1828), .C(n1620), .Y(n1629) );
  OAI21X1 U470 ( .A(n1036), .B(n984), .C(n1618), .Y(n1133) );
  NAND2X1 U471 ( .A(\mem<10><0> ), .B(n984), .Y(n1618) );
  OAI21X1 U472 ( .A(n1037), .B(n983), .C(n1617), .Y(n1132) );
  NAND2X1 U473 ( .A(\mem<10><1> ), .B(n984), .Y(n1617) );
  OAI21X1 U474 ( .A(n1038), .B(n983), .C(n1616), .Y(n1131) );
  NAND2X1 U475 ( .A(\mem<10><2> ), .B(n984), .Y(n1616) );
  OAI21X1 U476 ( .A(n1039), .B(n983), .C(n1615), .Y(n1130) );
  NAND2X1 U477 ( .A(\mem<10><3> ), .B(n984), .Y(n1615) );
  OAI21X1 U478 ( .A(n1040), .B(n983), .C(n1614), .Y(n1129) );
  NAND2X1 U479 ( .A(\mem<10><4> ), .B(n984), .Y(n1614) );
  OAI21X1 U480 ( .A(n1041), .B(n983), .C(n1613), .Y(n1128) );
  NAND2X1 U481 ( .A(\mem<10><5> ), .B(n984), .Y(n1613) );
  OAI21X1 U482 ( .A(n1042), .B(n983), .C(n1612), .Y(n1127) );
  NAND2X1 U483 ( .A(\mem<10><6> ), .B(n984), .Y(n1612) );
  OAI21X1 U484 ( .A(n1043), .B(n983), .C(n1611), .Y(n1126) );
  NAND2X1 U485 ( .A(\mem<10><7> ), .B(n984), .Y(n1611) );
  NAND3X1 U486 ( .A(n1766), .B(n1828), .C(n1651), .Y(n1619) );
  OAI21X1 U487 ( .A(n1028), .B(n982), .C(n1609), .Y(n1125) );
  NAND2X1 U488 ( .A(\mem<9><0> ), .B(n982), .Y(n1609) );
  OAI21X1 U489 ( .A(n1029), .B(n982), .C(n1608), .Y(n1124) );
  NAND2X1 U490 ( .A(\mem<9><1> ), .B(n982), .Y(n1608) );
  OAI21X1 U491 ( .A(n1030), .B(n982), .C(n1607), .Y(n1123) );
  NAND2X1 U492 ( .A(\mem<9><2> ), .B(n982), .Y(n1607) );
  OAI21X1 U493 ( .A(n1031), .B(n982), .C(n1606), .Y(n1122) );
  NAND2X1 U494 ( .A(\mem<9><3> ), .B(n982), .Y(n1606) );
  OAI21X1 U495 ( .A(n1032), .B(n982), .C(n1605), .Y(n1121) );
  NAND2X1 U496 ( .A(\mem<9><4> ), .B(n982), .Y(n1605) );
  OAI21X1 U497 ( .A(n1033), .B(n982), .C(n1604), .Y(n1120) );
  NAND2X1 U498 ( .A(\mem<9><5> ), .B(n982), .Y(n1604) );
  OAI21X1 U499 ( .A(n1034), .B(n982), .C(n1603), .Y(n1119) );
  NAND2X1 U500 ( .A(\mem<9><6> ), .B(n982), .Y(n1603) );
  OAI21X1 U501 ( .A(n1035), .B(n982), .C(n1602), .Y(n1118) );
  NAND2X1 U502 ( .A(\mem<9><7> ), .B(n982), .Y(n1602) );
  NAND3X1 U503 ( .A(n973), .B(n1828), .C(n1601), .Y(n1610) );
  OAI21X1 U504 ( .A(n1036), .B(n981), .C(n1599), .Y(n1117) );
  NAND2X1 U505 ( .A(\mem<8><0> ), .B(n981), .Y(n1599) );
  OAI21X1 U506 ( .A(n1037), .B(n980), .C(n1598), .Y(n1116) );
  NAND2X1 U507 ( .A(\mem<8><1> ), .B(n981), .Y(n1598) );
  OAI21X1 U508 ( .A(n1038), .B(n980), .C(n1597), .Y(n1115) );
  NAND2X1 U509 ( .A(\mem<8><2> ), .B(n981), .Y(n1597) );
  OAI21X1 U510 ( .A(n1039), .B(n980), .C(n1596), .Y(n1114) );
  NAND2X1 U511 ( .A(\mem<8><3> ), .B(n981), .Y(n1596) );
  OAI21X1 U512 ( .A(n1040), .B(n980), .C(n1595), .Y(n1113) );
  NAND2X1 U513 ( .A(\mem<8><4> ), .B(n981), .Y(n1595) );
  OAI21X1 U514 ( .A(n1041), .B(n980), .C(n1594), .Y(n1112) );
  NAND2X1 U515 ( .A(\mem<8><5> ), .B(n981), .Y(n1594) );
  OAI21X1 U516 ( .A(n1042), .B(n980), .C(n1593), .Y(n1111) );
  NAND2X1 U517 ( .A(\mem<8><6> ), .B(n981), .Y(n1593) );
  OAI21X1 U518 ( .A(n1043), .B(n980), .C(n1592), .Y(n1110) );
  NAND2X1 U519 ( .A(\mem<8><7> ), .B(n981), .Y(n1592) );
  NAND3X1 U520 ( .A(n1766), .B(n1828), .C(n1631), .Y(n1600) );
  OAI21X1 U521 ( .A(n1028), .B(n979), .C(n1589), .Y(n1109) );
  NAND2X1 U522 ( .A(\mem<7><0> ), .B(n979), .Y(n1589) );
  OAI21X1 U523 ( .A(n1029), .B(n979), .C(n1588), .Y(n1108) );
  NAND2X1 U524 ( .A(\mem<7><1> ), .B(n979), .Y(n1588) );
  OAI21X1 U525 ( .A(n1030), .B(n979), .C(n1587), .Y(n1107) );
  NAND2X1 U526 ( .A(\mem<7><2> ), .B(n979), .Y(n1587) );
  OAI21X1 U527 ( .A(n1031), .B(n979), .C(n1586), .Y(n1106) );
  NAND2X1 U528 ( .A(\mem<7><3> ), .B(n979), .Y(n1586) );
  OAI21X1 U529 ( .A(n1032), .B(n979), .C(n1585), .Y(n1105) );
  NAND2X1 U530 ( .A(\mem<7><4> ), .B(n979), .Y(n1585) );
  OAI21X1 U531 ( .A(n1033), .B(n979), .C(n1584), .Y(n1104) );
  NAND2X1 U532 ( .A(\mem<7><5> ), .B(n979), .Y(n1584) );
  OAI21X1 U533 ( .A(n1034), .B(n979), .C(n1583), .Y(n1103) );
  NAND2X1 U534 ( .A(\mem<7><6> ), .B(n979), .Y(n1583) );
  OAI21X1 U535 ( .A(n1035), .B(n979), .C(n1582), .Y(n1102) );
  NAND2X1 U536 ( .A(\mem<7><7> ), .B(n979), .Y(n1582) );
  NAND3X1 U537 ( .A(n973), .B(n1828), .C(n1581), .Y(n1590) );
  OAI21X1 U538 ( .A(n1036), .B(n978), .C(n1579), .Y(n1101) );
  NAND2X1 U539 ( .A(\mem<6><0> ), .B(n978), .Y(n1579) );
  OAI21X1 U540 ( .A(n1037), .B(n978), .C(n1578), .Y(n1100) );
  NAND2X1 U541 ( .A(\mem<6><1> ), .B(n978), .Y(n1578) );
  OAI21X1 U542 ( .A(n1038), .B(n978), .C(n1577), .Y(n1099) );
  NAND2X1 U543 ( .A(\mem<6><2> ), .B(n978), .Y(n1577) );
  OAI21X1 U544 ( .A(n1039), .B(n978), .C(n1576), .Y(n1098) );
  NAND2X1 U545 ( .A(\mem<6><3> ), .B(n978), .Y(n1576) );
  OAI21X1 U546 ( .A(n1040), .B(n978), .C(n1575), .Y(n1097) );
  NAND2X1 U547 ( .A(\mem<6><4> ), .B(n978), .Y(n1575) );
  OAI21X1 U548 ( .A(n1041), .B(n978), .C(n1574), .Y(n1096) );
  NAND2X1 U549 ( .A(\mem<6><5> ), .B(n978), .Y(n1574) );
  OAI21X1 U550 ( .A(n1042), .B(n978), .C(n1573), .Y(n1095) );
  NAND2X1 U551 ( .A(\mem<6><6> ), .B(n978), .Y(n1573) );
  OAI21X1 U552 ( .A(n1043), .B(n978), .C(n1572), .Y(n1094) );
  NAND2X1 U553 ( .A(\mem<6><7> ), .B(n978), .Y(n1572) );
  NAND3X1 U554 ( .A(n969), .B(n1828), .C(n1651), .Y(n1580) );
  OAI21X1 U555 ( .A(n1028), .B(n977), .C(n1570), .Y(n1093) );
  NAND2X1 U556 ( .A(\mem<5><0> ), .B(n977), .Y(n1570) );
  OAI21X1 U557 ( .A(n1029), .B(n977), .C(n1569), .Y(n1092) );
  NAND2X1 U558 ( .A(\mem<5><1> ), .B(n977), .Y(n1569) );
  OAI21X1 U559 ( .A(n1030), .B(n977), .C(n1568), .Y(n1091) );
  NAND2X1 U560 ( .A(\mem<5><2> ), .B(n977), .Y(n1568) );
  OAI21X1 U561 ( .A(n1031), .B(n977), .C(n1567), .Y(n1090) );
  NAND2X1 U562 ( .A(\mem<5><3> ), .B(n977), .Y(n1567) );
  OAI21X1 U563 ( .A(n1032), .B(n977), .C(n1566), .Y(n1089) );
  NAND2X1 U564 ( .A(\mem<5><4> ), .B(n977), .Y(n1566) );
  OAI21X1 U565 ( .A(n1033), .B(n977), .C(n1565), .Y(n1088) );
  NAND2X1 U566 ( .A(\mem<5><5> ), .B(n977), .Y(n1565) );
  OAI21X1 U567 ( .A(n1034), .B(n977), .C(n1564), .Y(n1087) );
  NAND2X1 U568 ( .A(\mem<5><6> ), .B(n977), .Y(n1564) );
  OAI21X1 U569 ( .A(n1035), .B(n977), .C(n1563), .Y(n1086) );
  NAND2X1 U570 ( .A(\mem<5><7> ), .B(n977), .Y(n1563) );
  NAND3X1 U571 ( .A(n973), .B(n1828), .C(n1562), .Y(n1571) );
  OAI21X1 U572 ( .A(n1036), .B(n976), .C(n1560), .Y(n1085) );
  NAND2X1 U573 ( .A(\mem<4><0> ), .B(n976), .Y(n1560) );
  OAI21X1 U574 ( .A(n1037), .B(n976), .C(n1559), .Y(n1084) );
  NAND2X1 U575 ( .A(\mem<4><1> ), .B(n976), .Y(n1559) );
  OAI21X1 U576 ( .A(n1038), .B(n976), .C(n1558), .Y(n1083) );
  NAND2X1 U577 ( .A(\mem<4><2> ), .B(n976), .Y(n1558) );
  OAI21X1 U578 ( .A(n1039), .B(n976), .C(n1557), .Y(n1082) );
  NAND2X1 U579 ( .A(\mem<4><3> ), .B(n976), .Y(n1557) );
  OAI21X1 U580 ( .A(n1040), .B(n976), .C(n1556), .Y(n1081) );
  NAND2X1 U581 ( .A(\mem<4><4> ), .B(n976), .Y(n1556) );
  OAI21X1 U582 ( .A(n1041), .B(n976), .C(n1555), .Y(n1080) );
  NAND2X1 U583 ( .A(\mem<4><5> ), .B(n976), .Y(n1555) );
  OAI21X1 U584 ( .A(n1042), .B(n976), .C(n1554), .Y(n1079) );
  NAND2X1 U585 ( .A(\mem<4><6> ), .B(n976), .Y(n1554) );
  OAI21X1 U586 ( .A(n1043), .B(n976), .C(n1553), .Y(n1078) );
  NAND2X1 U587 ( .A(\mem<4><7> ), .B(n976), .Y(n1553) );
  NAND3X1 U588 ( .A(n969), .B(n1828), .C(n1631), .Y(n1561) );
  OAI21X1 U590 ( .A(n1028), .B(n975), .C(n1550), .Y(n1077) );
  NAND2X1 U591 ( .A(\mem<3><0> ), .B(n975), .Y(n1550) );
  OAI21X1 U592 ( .A(n1029), .B(n975), .C(n1549), .Y(n1076) );
  NAND2X1 U593 ( .A(\mem<3><1> ), .B(n975), .Y(n1549) );
  OAI21X1 U594 ( .A(n1030), .B(n975), .C(n1548), .Y(n1075) );
  NAND2X1 U595 ( .A(\mem<3><2> ), .B(n975), .Y(n1548) );
  OAI21X1 U596 ( .A(n1031), .B(n975), .C(n1547), .Y(n1074) );
  NAND2X1 U597 ( .A(\mem<3><3> ), .B(n975), .Y(n1547) );
  OAI21X1 U598 ( .A(n1032), .B(n975), .C(n1546), .Y(n1073) );
  NAND2X1 U599 ( .A(\mem<3><4> ), .B(n975), .Y(n1546) );
  OAI21X1 U600 ( .A(n1033), .B(n975), .C(n1545), .Y(n1072) );
  NAND2X1 U601 ( .A(\mem<3><5> ), .B(n975), .Y(n1545) );
  OAI21X1 U602 ( .A(n1034), .B(n975), .C(n1544), .Y(n1071) );
  NAND2X1 U603 ( .A(\mem<3><6> ), .B(n975), .Y(n1544) );
  OAI21X1 U604 ( .A(n1035), .B(n975), .C(n1543), .Y(n1070) );
  NAND2X1 U605 ( .A(\mem<3><7> ), .B(n975), .Y(n1543) );
  NAND3X1 U606 ( .A(n973), .B(n1828), .C(n1542), .Y(n1551) );
  OAI21X1 U607 ( .A(n1036), .B(n974), .C(n1540), .Y(n1069) );
  NAND2X1 U608 ( .A(\mem<2><0> ), .B(n974), .Y(n1540) );
  OAI21X1 U609 ( .A(n1037), .B(n974), .C(n1539), .Y(n1068) );
  NAND2X1 U610 ( .A(\mem<2><1> ), .B(n974), .Y(n1539) );
  OAI21X1 U611 ( .A(n1038), .B(n974), .C(n1538), .Y(n1067) );
  NAND2X1 U612 ( .A(\mem<2><2> ), .B(n974), .Y(n1538) );
  OAI21X1 U613 ( .A(n1039), .B(n974), .C(n1537), .Y(n1066) );
  NAND2X1 U614 ( .A(\mem<2><3> ), .B(n974), .Y(n1537) );
  OAI21X1 U615 ( .A(n1040), .B(n974), .C(n1536), .Y(n1065) );
  NAND2X1 U616 ( .A(\mem<2><4> ), .B(n974), .Y(n1536) );
  OAI21X1 U617 ( .A(n1041), .B(n974), .C(n1535), .Y(n1064) );
  NAND2X1 U618 ( .A(\mem<2><5> ), .B(n974), .Y(n1535) );
  OAI21X1 U619 ( .A(n1042), .B(n974), .C(n1534), .Y(n1063) );
  NAND2X1 U620 ( .A(\mem<2><6> ), .B(n974), .Y(n1534) );
  OAI21X1 U621 ( .A(n1043), .B(n974), .C(n1533), .Y(n1062) );
  NAND2X1 U622 ( .A(\mem<2><7> ), .B(n974), .Y(n1533) );
  NAND3X1 U623 ( .A(n967), .B(n1828), .C(n1651), .Y(n1541) );
  OAI21X1 U624 ( .A(n1028), .B(n8), .C(n1532), .Y(n1061) );
  NAND2X1 U625 ( .A(\mem<1><0> ), .B(n8), .Y(n1532) );
  OAI21X1 U626 ( .A(n1029), .B(n8), .C(n1531), .Y(n1060) );
  NAND2X1 U627 ( .A(\mem<1><1> ), .B(n8), .Y(n1531) );
  OAI21X1 U628 ( .A(n1030), .B(n8), .C(n1530), .Y(n1059) );
  NAND2X1 U629 ( .A(\mem<1><2> ), .B(n8), .Y(n1530) );
  OAI21X1 U630 ( .A(n1031), .B(n8), .C(n1529), .Y(n1058) );
  NAND2X1 U631 ( .A(\mem<1><3> ), .B(n8), .Y(n1529) );
  OAI21X1 U632 ( .A(n1032), .B(n8), .C(n1528), .Y(n1057) );
  NAND2X1 U633 ( .A(\mem<1><4> ), .B(n8), .Y(n1528) );
  OAI21X1 U634 ( .A(n1033), .B(n8), .C(n1527), .Y(n1056) );
  NAND2X1 U635 ( .A(\mem<1><5> ), .B(n8), .Y(n1527) );
  OAI21X1 U636 ( .A(n1034), .B(n8), .C(n1526), .Y(n1055) );
  NAND2X1 U637 ( .A(\mem<1><6> ), .B(n8), .Y(n1526) );
  OAI21X1 U638 ( .A(n1035), .B(n8), .C(n1525), .Y(n1054) );
  NAND2X1 U639 ( .A(\mem<1><7> ), .B(n8), .Y(n1525) );
  NOR2X1 U641 ( .A(n965), .B(\addr_1c<4> ), .Y(n1818) );
  OAI21X1 U642 ( .A(n1036), .B(n972), .C(n1522), .Y(n1053) );
  NAND2X1 U643 ( .A(\mem<0><0> ), .B(n972), .Y(n1522) );
  OAI21X1 U644 ( .A(n1037), .B(n972), .C(n1521), .Y(n1052) );
  NAND2X1 U645 ( .A(\mem<0><1> ), .B(n972), .Y(n1521) );
  OAI21X1 U646 ( .A(n1038), .B(n972), .C(n1520), .Y(n1051) );
  NAND2X1 U647 ( .A(\mem<0><2> ), .B(n972), .Y(n1520) );
  OAI21X1 U648 ( .A(n1039), .B(n972), .C(n1519), .Y(n1050) );
  NAND2X1 U649 ( .A(\mem<0><3> ), .B(n972), .Y(n1519) );
  OAI21X1 U650 ( .A(n1040), .B(n972), .C(n1518), .Y(n1049) );
  NAND2X1 U651 ( .A(\mem<0><4> ), .B(n972), .Y(n1518) );
  OAI21X1 U652 ( .A(n1041), .B(n972), .C(n1517), .Y(n1048) );
  NAND2X1 U653 ( .A(\mem<0><5> ), .B(n972), .Y(n1517) );
  OAI21X1 U654 ( .A(n1042), .B(n972), .C(n1516), .Y(n1047) );
  NAND2X1 U655 ( .A(\mem<0><6> ), .B(n972), .Y(n1516) );
  OAI21X1 U656 ( .A(n1043), .B(n972), .C(n1515), .Y(n1046) );
  NAND2X1 U657 ( .A(\mem<0><7> ), .B(n972), .Y(n1515) );
  NAND3X1 U658 ( .A(n967), .B(n1828), .C(n1631), .Y(n1523) );
  NOR3X1 U661 ( .A(n1511), .B(\addr_1c<7> ), .C(\addr_1c<6> ), .Y(n1512) );
  NOR3X1 U662 ( .A(n1510), .B(\addr_1c<11> ), .C(\addr_1c<10> ), .Y(n1513) );
  AOI21X1 U663 ( .A(n461), .B(n1509), .C(n963), .Y(n1838) );
  OAI21X1 U665 ( .A(rd), .B(n1508), .C(wr), .Y(n1509) );
  NAND3X1 U667 ( .A(n1507), .B(n1023), .C(n1506), .Y(n1508) );
  NOR3X1 U668 ( .A(rd1), .B(rd3), .C(rd2), .Y(n1506) );
  NOR2X1 U669 ( .A(wr3), .B(wr2), .Y(n1507) );
  AOI21X1 U670 ( .A(n448), .B(n1504), .C(n1014), .Y(\data_out_1c<9> ) );
  NOR3X1 U671 ( .A(n2), .B(n1503), .C(n4), .Y(n1504) );
  AOI22X1 U673 ( .A(\mem<16><1> ), .B(n1786), .C(\mem<0><1> ), .D(n1631), .Y(
        n1501) );
  AOI22X1 U674 ( .A(\mem<18><1> ), .B(n1806), .C(\mem<2><1> ), .D(n1651), .Y(
        n1502) );
  AOI22X1 U676 ( .A(\mem<20><1> ), .B(n1786), .C(\mem<4><1> ), .D(n1631), .Y(
        n1499) );
  AOI22X1 U677 ( .A(\mem<22><1> ), .B(n1806), .C(\mem<6><1> ), .D(n1651), .Y(
        n1500) );
  AOI22X1 U678 ( .A(n1591), .B(n892), .C(n1630), .D(n932), .Y(n1505) );
  AOI22X1 U680 ( .A(\mem<28><1> ), .B(n1786), .C(\mem<12><1> ), .D(n1631), .Y(
        n1497) );
  AOI22X1 U681 ( .A(\mem<30><1> ), .B(n1806), .C(\mem<14><1> ), .D(n1651), .Y(
        n1498) );
  AOI22X1 U683 ( .A(\mem<24><1> ), .B(n1786), .C(\mem<8><1> ), .D(n1631), .Y(
        n1495) );
  AOI22X1 U684 ( .A(\mem<26><1> ), .B(n1806), .C(\mem<10><1> ), .D(n1651), .Y(
        n1496) );
  AOI21X1 U685 ( .A(n447), .B(n1493), .C(n1014), .Y(\data_out_1c<8> ) );
  NOR3X1 U686 ( .A(n939), .B(n1491), .C(n950), .Y(n1493) );
  AOI21X1 U687 ( .A(n1489), .B(n1488), .C(n971), .Y(n1490) );
  AOI22X1 U688 ( .A(\mem<16><0> ), .B(n1786), .C(\mem<0><0> ), .D(n1631), .Y(
        n1488) );
  AOI22X1 U689 ( .A(\mem<18><0> ), .B(n1806), .C(\mem<2><0> ), .D(n1651), .Y(
        n1489) );
  AOI21X1 U690 ( .A(n1487), .B(n1486), .C(n970), .Y(n1492) );
  AOI22X1 U691 ( .A(\mem<20><0> ), .B(n1786), .C(\mem<4><0> ), .D(n1631), .Y(
        n1486) );
  AOI22X1 U692 ( .A(\mem<22><0> ), .B(n1806), .C(\mem<6><0> ), .D(n1651), .Y(
        n1487) );
  AOI22X1 U693 ( .A(n1591), .B(n890), .C(n1630), .D(n930), .Y(n1494) );
  AOI22X1 U695 ( .A(\mem<28><0> ), .B(n1786), .C(\mem<12><0> ), .D(n1631), .Y(
        n1484) );
  AOI22X1 U696 ( .A(\mem<30><0> ), .B(n1806), .C(\mem<14><0> ), .D(n1651), .Y(
        n1485) );
  AOI22X1 U698 ( .A(\mem<24><0> ), .B(n1786), .C(\mem<8><0> ), .D(n1631), .Y(
        n1482) );
  AOI22X1 U699 ( .A(\mem<26><0> ), .B(n1806), .C(\mem<10><0> ), .D(n1651), .Y(
        n1483) );
  OAI21X1 U700 ( .A(n23), .B(n50), .C(rd1), .Y(n1481) );
  AOI22X1 U702 ( .A(\mem<17><7> ), .B(n1680), .C(\mem<19><7> ), .D(n1699), .Y(
        n1476) );
  AOI22X1 U703 ( .A(\mem<21><7> ), .B(n1718), .C(\mem<23><7> ), .D(n1737), .Y(
        n1477) );
  AOI22X1 U704 ( .A(\mem<25><7> ), .B(n1756), .C(\mem<27><7> ), .D(n1776), .Y(
        n1479) );
  AOI22X1 U705 ( .A(\mem<29><7> ), .B(n1796), .C(\mem<31><7> ), .D(n1817), .Y(
        n1480) );
  AOI22X1 U707 ( .A(\mem<1><7> ), .B(n1524), .C(\mem<3><7> ), .D(n1542), .Y(
        n1471) );
  AOI22X1 U708 ( .A(\mem<5><7> ), .B(n1562), .C(\mem<7><7> ), .D(n1581), .Y(
        n1472) );
  AOI22X1 U709 ( .A(\mem<9><7> ), .B(n1601), .C(\mem<11><7> ), .D(n1620), .Y(
        n1474) );
  AOI22X1 U710 ( .A(\mem<13><7> ), .B(n1641), .C(\mem<15><7> ), .D(n1661), .Y(
        n1475) );
  OAI21X1 U711 ( .A(n21), .B(n37), .C(rd1), .Y(n1470) );
  AOI22X1 U713 ( .A(\mem<17><6> ), .B(n1680), .C(\mem<19><6> ), .D(n1699), .Y(
        n1465) );
  AOI22X1 U714 ( .A(\mem<21><6> ), .B(n1718), .C(\mem<23><6> ), .D(n1737), .Y(
        n1466) );
  AOI22X1 U715 ( .A(\mem<25><6> ), .B(n1756), .C(\mem<27><6> ), .D(n1776), .Y(
        n1468) );
  AOI22X1 U716 ( .A(\mem<29><6> ), .B(n1796), .C(\mem<31><6> ), .D(n1817), .Y(
        n1469) );
  AOI22X1 U718 ( .A(\mem<1><6> ), .B(n1524), .C(\mem<3><6> ), .D(n1542), .Y(
        n1460) );
  AOI22X1 U719 ( .A(\mem<5><6> ), .B(n1562), .C(\mem<7><6> ), .D(n1581), .Y(
        n1461) );
  AOI22X1 U720 ( .A(\mem<9><6> ), .B(n1601), .C(\mem<11><6> ), .D(n1620), .Y(
        n1463) );
  AOI22X1 U721 ( .A(\mem<13><6> ), .B(n1641), .C(\mem<15><6> ), .D(n1661), .Y(
        n1464) );
  OAI21X1 U722 ( .A(n19), .B(n35), .C(rd1), .Y(n1459) );
  AOI22X1 U724 ( .A(\mem<17><5> ), .B(n1680), .C(\mem<19><5> ), .D(n1699), .Y(
        n1454) );
  AOI22X1 U725 ( .A(\mem<21><5> ), .B(n1718), .C(\mem<23><5> ), .D(n1737), .Y(
        n1455) );
  AOI22X1 U726 ( .A(\mem<25><5> ), .B(n1756), .C(\mem<27><5> ), .D(n1776), .Y(
        n1457) );
  AOI22X1 U727 ( .A(\mem<29><5> ), .B(n1796), .C(\mem<31><5> ), .D(n1817), .Y(
        n1458) );
  AOI22X1 U729 ( .A(\mem<1><5> ), .B(n1524), .C(\mem<3><5> ), .D(n1542), .Y(
        n1449) );
  AOI22X1 U730 ( .A(\mem<5><5> ), .B(n1562), .C(\mem<7><5> ), .D(n1581), .Y(
        n1450) );
  AOI22X1 U731 ( .A(\mem<9><5> ), .B(n1601), .C(\mem<11><5> ), .D(n1620), .Y(
        n1452) );
  AOI22X1 U732 ( .A(\mem<13><5> ), .B(n1641), .C(\mem<15><5> ), .D(n1661), .Y(
        n1453) );
  OAI21X1 U733 ( .A(n17), .B(n33), .C(rd1), .Y(n1448) );
  AOI22X1 U735 ( .A(\mem<17><4> ), .B(n1680), .C(\mem<19><4> ), .D(n1699), .Y(
        n1443) );
  AOI22X1 U736 ( .A(\mem<21><4> ), .B(n1718), .C(\mem<23><4> ), .D(n1737), .Y(
        n1444) );
  AOI22X1 U737 ( .A(\mem<25><4> ), .B(n1756), .C(\mem<27><4> ), .D(n1776), .Y(
        n1446) );
  AOI22X1 U738 ( .A(\mem<29><4> ), .B(n1796), .C(\mem<31><4> ), .D(n1817), .Y(
        n1447) );
  AOI22X1 U740 ( .A(\mem<1><4> ), .B(n1524), .C(\mem<3><4> ), .D(n1542), .Y(
        n1438) );
  AOI22X1 U741 ( .A(\mem<5><4> ), .B(n1562), .C(\mem<7><4> ), .D(n1581), .Y(
        n1439) );
  AOI22X1 U742 ( .A(\mem<9><4> ), .B(n1601), .C(\mem<11><4> ), .D(n1620), .Y(
        n1441) );
  AOI22X1 U743 ( .A(\mem<13><4> ), .B(n1641), .C(\mem<15><4> ), .D(n1661), .Y(
        n1442) );
  OAI21X1 U744 ( .A(n15), .B(n31), .C(rd1), .Y(n1437) );
  AOI22X1 U746 ( .A(\mem<17><3> ), .B(n1680), .C(\mem<19><3> ), .D(n1699), .Y(
        n1432) );
  AOI22X1 U747 ( .A(\mem<21><3> ), .B(n1718), .C(\mem<23><3> ), .D(n1737), .Y(
        n1433) );
  AOI22X1 U748 ( .A(\mem<25><3> ), .B(n1756), .C(\mem<27><3> ), .D(n1776), .Y(
        n1435) );
  AOI22X1 U749 ( .A(\mem<29><3> ), .B(n1796), .C(\mem<31><3> ), .D(n1817), .Y(
        n1436) );
  AOI22X1 U751 ( .A(\mem<1><3> ), .B(n1524), .C(\mem<3><3> ), .D(n1542), .Y(
        n1427) );
  AOI22X1 U752 ( .A(\mem<5><3> ), .B(n1562), .C(\mem<7><3> ), .D(n1581), .Y(
        n1428) );
  AOI22X1 U753 ( .A(\mem<9><3> ), .B(n1601), .C(\mem<11><3> ), .D(n1620), .Y(
        n1430) );
  AOI22X1 U754 ( .A(\mem<13><3> ), .B(n1641), .C(\mem<15><3> ), .D(n1661), .Y(
        n1431) );
  OAI21X1 U755 ( .A(n13), .B(n29), .C(rd1), .Y(n1426) );
  AOI22X1 U757 ( .A(\mem<17><2> ), .B(n1680), .C(\mem<19><2> ), .D(n1699), .Y(
        n1421) );
  AOI22X1 U758 ( .A(\mem<21><2> ), .B(n1718), .C(\mem<23><2> ), .D(n1737), .Y(
        n1422) );
  AOI22X1 U759 ( .A(\mem<25><2> ), .B(n1756), .C(\mem<27><2> ), .D(n1776), .Y(
        n1424) );
  AOI22X1 U760 ( .A(\mem<29><2> ), .B(n1796), .C(\mem<31><2> ), .D(n1817), .Y(
        n1425) );
  AOI22X1 U762 ( .A(\mem<1><2> ), .B(n1524), .C(\mem<3><2> ), .D(n1542), .Y(
        n1416) );
  AOI22X1 U763 ( .A(\mem<5><2> ), .B(n1562), .C(\mem<7><2> ), .D(n1581), .Y(
        n1417) );
  AOI22X1 U764 ( .A(\mem<9><2> ), .B(n1601), .C(\mem<11><2> ), .D(n1620), .Y(
        n1419) );
  AOI22X1 U765 ( .A(\mem<13><2> ), .B(n1641), .C(\mem<15><2> ), .D(n1661), .Y(
        n1420) );
  OAI21X1 U766 ( .A(n11), .B(n27), .C(rd1), .Y(n1415) );
  AOI22X1 U768 ( .A(\mem<17><1> ), .B(n1680), .C(\mem<19><1> ), .D(n1699), .Y(
        n1410) );
  AOI22X1 U769 ( .A(\mem<21><1> ), .B(n1718), .C(\mem<23><1> ), .D(n1737), .Y(
        n1411) );
  AOI22X1 U770 ( .A(\mem<25><1> ), .B(n1756), .C(\mem<27><1> ), .D(n1776), .Y(
        n1413) );
  AOI22X1 U771 ( .A(\mem<29><1> ), .B(n1796), .C(\mem<31><1> ), .D(n1817), .Y(
        n1414) );
  AOI22X1 U773 ( .A(\mem<1><1> ), .B(n1524), .C(\mem<3><1> ), .D(n1542), .Y(
        n1405) );
  AOI22X1 U774 ( .A(\mem<5><1> ), .B(n1562), .C(\mem<7><1> ), .D(n1581), .Y(
        n1406) );
  AOI22X1 U775 ( .A(\mem<9><1> ), .B(n1601), .C(\mem<11><1> ), .D(n1620), .Y(
        n1408) );
  AOI22X1 U776 ( .A(\mem<13><1> ), .B(n1641), .C(\mem<15><1> ), .D(n1661), .Y(
        n1409) );
  AOI21X1 U777 ( .A(n435), .B(n1403), .C(n1014), .Y(\data_out_1c<15> ) );
  NOR3X1 U778 ( .A(n938), .B(n1401), .C(n949), .Y(n1403) );
  AOI21X1 U779 ( .A(n1399), .B(n1398), .C(n971), .Y(n1400) );
  AOI22X1 U780 ( .A(\mem<16><7> ), .B(n1786), .C(\mem<0><7> ), .D(n1631), .Y(
        n1398) );
  AOI22X1 U781 ( .A(\mem<18><7> ), .B(n1806), .C(\mem<2><7> ), .D(n1651), .Y(
        n1399) );
  AOI21X1 U782 ( .A(n1397), .B(n1396), .C(n970), .Y(n1402) );
  AOI22X1 U783 ( .A(\mem<20><7> ), .B(n1786), .C(\mem<4><7> ), .D(n1631), .Y(
        n1396) );
  AOI22X1 U784 ( .A(\mem<22><7> ), .B(n1806), .C(\mem<6><7> ), .D(n1651), .Y(
        n1397) );
  AOI22X1 U785 ( .A(n1591), .B(n888), .C(n1630), .D(n928), .Y(n1404) );
  AOI22X1 U787 ( .A(\mem<28><7> ), .B(n1786), .C(\mem<12><7> ), .D(n1631), .Y(
        n1394) );
  AOI22X1 U788 ( .A(\mem<30><7> ), .B(n1806), .C(\mem<14><7> ), .D(n1651), .Y(
        n1395) );
  AOI22X1 U790 ( .A(\mem<24><7> ), .B(n1786), .C(\mem<8><7> ), .D(n1631), .Y(
        n1392) );
  AOI22X1 U791 ( .A(\mem<26><7> ), .B(n1806), .C(\mem<10><7> ), .D(n1651), .Y(
        n1393) );
  AOI21X1 U792 ( .A(n434), .B(n1390), .C(n1014), .Y(\data_out_1c<14> ) );
  NOR3X1 U793 ( .A(n937), .B(n1388), .C(n948), .Y(n1390) );
  AOI21X1 U794 ( .A(n1386), .B(n1385), .C(n971), .Y(n1387) );
  AOI22X1 U795 ( .A(\mem<16><6> ), .B(n1786), .C(\mem<0><6> ), .D(n1631), .Y(
        n1385) );
  AOI22X1 U796 ( .A(\mem<18><6> ), .B(n1806), .C(\mem<2><6> ), .D(n1651), .Y(
        n1386) );
  AOI21X1 U797 ( .A(n1384), .B(n1383), .C(n970), .Y(n1389) );
  AOI22X1 U798 ( .A(\mem<20><6> ), .B(n1786), .C(\mem<4><6> ), .D(n1631), .Y(
        n1383) );
  AOI22X1 U799 ( .A(\mem<22><6> ), .B(n1806), .C(\mem<6><6> ), .D(n1651), .Y(
        n1384) );
  AOI22X1 U800 ( .A(n1591), .B(n886), .C(n1630), .D(n926), .Y(n1391) );
  AOI22X1 U802 ( .A(\mem<28><6> ), .B(n1786), .C(\mem<12><6> ), .D(n1631), .Y(
        n1381) );
  AOI22X1 U803 ( .A(\mem<30><6> ), .B(n1806), .C(\mem<14><6> ), .D(n1651), .Y(
        n1382) );
  AOI22X1 U805 ( .A(\mem<24><6> ), .B(n1786), .C(\mem<8><6> ), .D(n1631), .Y(
        n1379) );
  AOI22X1 U806 ( .A(\mem<26><6> ), .B(n1806), .C(\mem<10><6> ), .D(n1651), .Y(
        n1380) );
  AOI21X1 U807 ( .A(n422), .B(n1377), .C(n1014), .Y(\data_out_1c<13> ) );
  NOR3X1 U808 ( .A(n936), .B(n1375), .C(n947), .Y(n1377) );
  AOI21X1 U809 ( .A(n1373), .B(n1372), .C(n971), .Y(n1374) );
  AOI22X1 U810 ( .A(\mem<16><5> ), .B(n1786), .C(\mem<0><5> ), .D(n1631), .Y(
        n1372) );
  AOI22X1 U811 ( .A(\mem<18><5> ), .B(n1806), .C(\mem<2><5> ), .D(n1651), .Y(
        n1373) );
  AOI21X1 U812 ( .A(n1371), .B(n1370), .C(n970), .Y(n1376) );
  AOI22X1 U813 ( .A(\mem<20><5> ), .B(n1786), .C(\mem<4><5> ), .D(n1631), .Y(
        n1370) );
  AOI22X1 U814 ( .A(\mem<22><5> ), .B(n1806), .C(\mem<6><5> ), .D(n1651), .Y(
        n1371) );
  AOI22X1 U815 ( .A(n1591), .B(n884), .C(n1630), .D(n924), .Y(n1378) );
  AOI22X1 U817 ( .A(\mem<28><5> ), .B(n1786), .C(\mem<12><5> ), .D(n1631), .Y(
        n1368) );
  AOI22X1 U818 ( .A(\mem<30><5> ), .B(n1806), .C(\mem<14><5> ), .D(n1651), .Y(
        n1369) );
  AOI22X1 U820 ( .A(\mem<24><5> ), .B(n1786), .C(\mem<8><5> ), .D(n1631), .Y(
        n1366) );
  AOI22X1 U821 ( .A(\mem<26><5> ), .B(n1806), .C(\mem<10><5> ), .D(n1651), .Y(
        n1367) );
  AOI21X1 U822 ( .A(n421), .B(n1364), .C(n1014), .Y(\data_out_1c<12> ) );
  NOR3X1 U823 ( .A(n935), .B(n1362), .C(n946), .Y(n1364) );
  AOI21X1 U824 ( .A(n1360), .B(n1359), .C(n971), .Y(n1361) );
  AOI22X1 U825 ( .A(\mem<16><4> ), .B(n1786), .C(\mem<0><4> ), .D(n1631), .Y(
        n1359) );
  AOI22X1 U826 ( .A(\mem<18><4> ), .B(n1806), .C(\mem<2><4> ), .D(n1651), .Y(
        n1360) );
  AOI21X1 U827 ( .A(n1358), .B(n1357), .C(n970), .Y(n1363) );
  AOI22X1 U828 ( .A(\mem<20><4> ), .B(n1786), .C(\mem<4><4> ), .D(n1631), .Y(
        n1357) );
  AOI22X1 U829 ( .A(\mem<22><4> ), .B(n1806), .C(\mem<6><4> ), .D(n1651), .Y(
        n1358) );
  AOI22X1 U830 ( .A(n1591), .B(n882), .C(n1630), .D(n922), .Y(n1365) );
  AOI22X1 U832 ( .A(\mem<28><4> ), .B(n1786), .C(\mem<12><4> ), .D(n1631), .Y(
        n1355) );
  AOI22X1 U833 ( .A(\mem<30><4> ), .B(n1806), .C(\mem<14><4> ), .D(n1651), .Y(
        n1356) );
  AOI22X1 U835 ( .A(\mem<24><4> ), .B(n1786), .C(\mem<8><4> ), .D(n1631), .Y(
        n1353) );
  AOI22X1 U836 ( .A(\mem<26><4> ), .B(n1806), .C(\mem<10><4> ), .D(n1651), .Y(
        n1354) );
  AOI21X1 U837 ( .A(n409), .B(n1351), .C(n1014), .Y(\data_out_1c<11> ) );
  NOR3X1 U838 ( .A(n934), .B(n1349), .C(n945), .Y(n1351) );
  AOI21X1 U839 ( .A(n1347), .B(n1346), .C(n971), .Y(n1348) );
  AOI22X1 U840 ( .A(\mem<16><3> ), .B(n1786), .C(\mem<0><3> ), .D(n1631), .Y(
        n1346) );
  AOI22X1 U841 ( .A(\mem<18><3> ), .B(n1806), .C(\mem<2><3> ), .D(n1651), .Y(
        n1347) );
  AOI21X1 U842 ( .A(n1345), .B(n1344), .C(n970), .Y(n1350) );
  AOI22X1 U843 ( .A(\mem<20><3> ), .B(n1786), .C(\mem<4><3> ), .D(n1631), .Y(
        n1344) );
  AOI22X1 U844 ( .A(\mem<22><3> ), .B(n1806), .C(\mem<6><3> ), .D(n1651), .Y(
        n1345) );
  AOI22X1 U845 ( .A(n1591), .B(n880), .C(n1630), .D(n920), .Y(n1352) );
  AOI22X1 U847 ( .A(\mem<28><3> ), .B(n1786), .C(\mem<12><3> ), .D(n1631), .Y(
        n1342) );
  AOI22X1 U848 ( .A(\mem<30><3> ), .B(n1806), .C(\mem<14><3> ), .D(n1651), .Y(
        n1343) );
  AOI22X1 U850 ( .A(\mem<24><3> ), .B(n1786), .C(\mem<8><3> ), .D(n1631), .Y(
        n1340) );
  AOI22X1 U851 ( .A(\mem<26><3> ), .B(n1806), .C(\mem<10><3> ), .D(n1651), .Y(
        n1341) );
  AOI21X1 U852 ( .A(n408), .B(n1338), .C(n1014), .Y(\data_out_1c<10> ) );
  NOR3X1 U853 ( .A(n933), .B(n1336), .C(n944), .Y(n1338) );
  AOI21X1 U854 ( .A(n1334), .B(n1333), .C(n971), .Y(n1335) );
  AOI22X1 U855 ( .A(\mem<16><2> ), .B(n1786), .C(\mem<0><2> ), .D(n1631), .Y(
        n1333) );
  AOI22X1 U856 ( .A(\mem<18><2> ), .B(n1806), .C(\mem<2><2> ), .D(n1651), .Y(
        n1334) );
  AOI21X1 U857 ( .A(n1332), .B(n1331), .C(n970), .Y(n1337) );
  AOI22X1 U858 ( .A(\mem<20><2> ), .B(n1786), .C(\mem<4><2> ), .D(n1631), .Y(
        n1331) );
  AOI22X1 U859 ( .A(\mem<22><2> ), .B(n1806), .C(\mem<6><2> ), .D(n1651), .Y(
        n1332) );
  AOI22X1 U860 ( .A(n1591), .B(n878), .C(n1630), .D(n918), .Y(n1339) );
  AOI22X1 U862 ( .A(\mem<28><2> ), .B(n1786), .C(\mem<12><2> ), .D(n1631), .Y(
        n1329) );
  AOI22X1 U863 ( .A(\mem<30><2> ), .B(n1806), .C(\mem<14><2> ), .D(n1651), .Y(
        n1330) );
  AOI22X1 U865 ( .A(\mem<24><2> ), .B(n1786), .C(\mem<8><2> ), .D(n1631), .Y(
        n1327) );
  AOI22X1 U866 ( .A(\mem<26><2> ), .B(n1806), .C(\mem<10><2> ), .D(n1651), .Y(
        n1328) );
  NOR2X1 U867 ( .A(\addr_1c<3> ), .B(\addr_1c<4> ), .Y(n1326) );
  NOR2X1 U868 ( .A(n1027), .B(\addr_1c<4> ), .Y(n1325) );
  OAI21X1 U869 ( .A(n9), .B(n25), .C(rd1), .Y(n1324) );
  AOI22X1 U871 ( .A(\mem<17><0> ), .B(n1680), .C(\mem<19><0> ), .D(n1699), .Y(
        n1319) );
  AOI22X1 U872 ( .A(\mem<21><0> ), .B(n1718), .C(\mem<23><0> ), .D(n1737), .Y(
        n1320) );
  AOI22X1 U873 ( .A(\mem<25><0> ), .B(n1756), .C(\mem<27><0> ), .D(n1776), .Y(
        n1322) );
  AOI22X1 U874 ( .A(\mem<29><0> ), .B(n1796), .C(\mem<31><0> ), .D(n1817), .Y(
        n1323) );
  AOI22X1 U876 ( .A(\mem<1><0> ), .B(n1524), .C(\mem<3><0> ), .D(n1542), .Y(
        n1312) );
  NAND2X1 U877 ( .A(n1025), .B(n1026), .Y(n1514) );
  AOI22X1 U878 ( .A(\mem<5><0> ), .B(n1562), .C(\mem<7><0> ), .D(n1581), .Y(
        n1313) );
  NAND2X1 U879 ( .A(\addr_1c<1> ), .B(n1026), .Y(n1552) );
  AOI22X1 U880 ( .A(\mem<9><0> ), .B(n1601), .C(\mem<11><0> ), .D(n1620), .Y(
        n1315) );
  AOI22X1 U881 ( .A(\mem<13><0> ), .B(n1641), .C(\mem<15><0> ), .D(n1661), .Y(
        n1316) );
  dff_54 ff0 ( .q(rd1), .d(rd0), .clk(clk), .rst(n1012) );
  dff_53 ff1 ( .q(wr1), .d(wr0), .clk(clk), .rst(n1012) );
  dff_52 \reg0[0]  ( .q(\addr_1c<0> ), .d(\addr<0> ), .clk(clk), .rst(n1012)
         );
  dff_51 \reg0[1]  ( .q(\addr_1c<1> ), .d(\addr<1> ), .clk(clk), .rst(n1012)
         );
  dff_50 \reg0[2]  ( .q(\addr_1c<2> ), .d(\addr<2> ), .clk(clk), .rst(n1012)
         );
  dff_49 \reg0[3]  ( .q(\addr_1c<3> ), .d(\addr<3> ), .clk(clk), .rst(n1012)
         );
  dff_48 \reg0[4]  ( .q(\addr_1c<4> ), .d(\addr<4> ), .clk(clk), .rst(n1012)
         );
  dff_47 \reg0[5]  ( .q(\addr_1c<5> ), .d(\addr<5> ), .clk(clk), .rst(n1012)
         );
  dff_46 \reg0[6]  ( .q(\addr_1c<6> ), .d(\addr<6> ), .clk(clk), .rst(n1012)
         );
  dff_45 \reg0[7]  ( .q(\addr_1c<7> ), .d(\addr<7> ), .clk(clk), .rst(n1012)
         );
  dff_44 \reg0[8]  ( .q(\addr_1c<8> ), .d(\addr<8> ), .clk(clk), .rst(n1012)
         );
  dff_43 \reg0[9]  ( .q(\addr_1c<9> ), .d(\addr<9> ), .clk(clk), .rst(n1012)
         );
  dff_42 \reg0[10]  ( .q(\addr_1c<10> ), .d(\addr<10> ), .clk(clk), .rst(n1012) );
  dff_41 \reg0[11]  ( .q(\addr_1c<11> ), .d(\addr<11> ), .clk(clk), .rst(n1012) );
  dff_40 \reg0[12]  ( .q(\addr_1c<12> ), .d(\addr<12> ), .clk(clk), .rst(n1012) );
  dff_39 \reg1[0]  ( .q(\data_in_1c<0> ), .d(\data_in<0> ), .clk(clk), .rst(
        n1012) );
  dff_38 \reg1[1]  ( .q(\data_in_1c<1> ), .d(\data_in<1> ), .clk(clk), .rst(
        n1012) );
  dff_37 \reg1[2]  ( .q(\data_in_1c<2> ), .d(\data_in<2> ), .clk(clk), .rst(
        n1012) );
  dff_36 \reg1[3]  ( .q(\data_in_1c<3> ), .d(\data_in<3> ), .clk(clk), .rst(
        n1012) );
  dff_35 \reg1[4]  ( .q(\data_in_1c<4> ), .d(\data_in<4> ), .clk(clk), .rst(
        n1012) );
  dff_34 \reg1[5]  ( .q(\data_in_1c<5> ), .d(\data_in<5> ), .clk(clk), .rst(
        n1012) );
  dff_33 \reg1[6]  ( .q(\data_in_1c<6> ), .d(\data_in<6> ), .clk(clk), .rst(
        n1012) );
  dff_32 \reg1[7]  ( .q(\data_in_1c<7> ), .d(\data_in<7> ), .clk(clk), .rst(
        n1012) );
  dff_31 \reg1[8]  ( .q(\data_in_1c<8> ), .d(\data_in<8> ), .clk(clk), .rst(
        n1012) );
  dff_30 \reg1[9]  ( .q(\data_in_1c<9> ), .d(\data_in<9> ), .clk(clk), .rst(
        n1012) );
  dff_29 \reg1[10]  ( .q(\data_in_1c<10> ), .d(\data_in<10> ), .clk(clk), 
        .rst(n1012) );
  dff_28 \reg1[11]  ( .q(\data_in_1c<11> ), .d(\data_in<11> ), .clk(clk), 
        .rst(n1012) );
  dff_27 \reg1[12]  ( .q(\data_in_1c<12> ), .d(\data_in<12> ), .clk(clk), 
        .rst(n1012) );
  dff_26 \reg1[13]  ( .q(\data_in_1c<13> ), .d(\data_in<13> ), .clk(clk), 
        .rst(n1012) );
  dff_25 \reg1[14]  ( .q(\data_in_1c<14> ), .d(\data_in<14> ), .clk(clk), 
        .rst(n1012) );
  dff_24 \reg1[15]  ( .q(\data_in_1c<15> ), .d(\data_in<15> ), .clk(clk), 
        .rst(n1012) );
  dff_23 \reg2[0]  ( .q(\data_out<0> ), .d(n1022), .clk(clk), .rst(n1012) );
  dff_22 \reg2[1]  ( .q(\data_out<1> ), .d(n1021), .clk(clk), .rst(n1012) );
  dff_21 \reg2[2]  ( .q(\data_out<2> ), .d(n1020), .clk(clk), .rst(n1012) );
  dff_20 \reg2[3]  ( .q(\data_out<3> ), .d(n1019), .clk(clk), .rst(n1012) );
  dff_19 \reg2[4]  ( .q(\data_out<4> ), .d(n1018), .clk(clk), .rst(n1012) );
  dff_18 \reg2[5]  ( .q(\data_out<5> ), .d(n1017), .clk(clk), .rst(n1012) );
  dff_17 \reg2[6]  ( .q(\data_out<6> ), .d(n1016), .clk(clk), .rst(n1012) );
  dff_16 \reg2[7]  ( .q(\data_out<7> ), .d(n1015), .clk(clk), .rst(n1012) );
  dff_15 \reg2[8]  ( .q(\data_out<8> ), .d(\data_out_1c<8> ), .clk(clk), .rst(
        n1012) );
  dff_14 \reg2[9]  ( .q(\data_out<9> ), .d(\data_out_1c<9> ), .clk(clk), .rst(
        n1012) );
  dff_13 \reg2[10]  ( .q(\data_out<10> ), .d(\data_out_1c<10> ), .clk(clk), 
        .rst(n1012) );
  dff_12 \reg2[11]  ( .q(\data_out<11> ), .d(\data_out_1c<11> ), .clk(clk), 
        .rst(n1012) );
  dff_11 \reg2[12]  ( .q(\data_out<12> ), .d(\data_out_1c<12> ), .clk(clk), 
        .rst(n1012) );
  dff_10 \reg2[13]  ( .q(\data_out<13> ), .d(\data_out_1c<13> ), .clk(clk), 
        .rst(n1012) );
  dff_9 \reg2[14]  ( .q(\data_out<14> ), .d(\data_out_1c<14> ), .clk(clk), 
        .rst(n1012) );
  dff_8 \reg2[15]  ( .q(\data_out<15> ), .d(\data_out_1c<15> ), .clk(clk), 
        .rst(n1012) );
  dff_7 ff2 ( .q(rd2), .d(rd1), .clk(clk), .rst(n1012) );
  dff_6 ff3 ( .q(wr2), .d(wr1), .clk(clk), .rst(n1012) );
  dff_5 ff4 ( .q(rd3), .d(rd2), .clk(clk), .rst(n1012) );
  dff_4 ff5 ( .q(wr3), .d(wr2), .clk(clk), .rst(n1012) );
  INVX1 U2 ( .A(rd), .Y(n1045) );
  OR2X1 U3 ( .A(\addr_1c<5> ), .B(\addr_1c<12> ), .Y(n1510) );
  AND2X1 U4 ( .A(\addr_1c<4> ), .B(n1524), .Y(n1827) );
  INVX1 U5 ( .A(\addr_1c<3> ), .Y(n1027) );
  INVX1 U6 ( .A(\addr_1c<2> ), .Y(n1026) );
  INVX1 U7 ( .A(wr1), .Y(n1023) );
  INVX1 U8 ( .A(\addr_1c<1> ), .Y(n1025) );
  OR2X1 U23 ( .A(\addr_1c<9> ), .B(\addr_1c<8> ), .Y(n1511) );
  AND2X1 U24 ( .A(\addr_1c<3> ), .B(\addr_1c<0> ), .Y(n1318) );
  AND2X1 U25 ( .A(\addr_1c<3> ), .B(n1024), .Y(n1317) );
  AND2X1 U26 ( .A(n1630), .B(n964), .Y(n1807) );
  AND2X1 U27 ( .A(n1591), .B(n964), .Y(n1766) );
  AND2X1 U28 ( .A(\addr_1c<0> ), .B(n1027), .Y(n1311) );
  AND2X1 U29 ( .A(n1024), .B(n1027), .Y(n1310) );
  INVX1 U35 ( .A(\addr_1c<0> ), .Y(n1024) );
  AND2X1 U36 ( .A(\addr_1c<2> ), .B(n1025), .Y(n1591) );
  AND2X1 U37 ( .A(\addr_1c<2> ), .B(\addr_1c<1> ), .Y(n1630) );
  AND2X1 U38 ( .A(n1317), .B(n1630), .Y(n1796) );
  AND2X1 U39 ( .A(n1591), .B(n1318), .Y(n1776) );
  AND2X1 U40 ( .A(n1591), .B(n1317), .Y(n1756) );
  AND2X1 U41 ( .A(n940), .B(n1318), .Y(n1737) );
  AND2X1 U42 ( .A(n940), .B(n1317), .Y(n1718) );
  AND2X1 U43 ( .A(n1318), .B(n951), .Y(n1699) );
  AND2X1 U44 ( .A(n1317), .B(n951), .Y(n1680) );
  AND2X1 U46 ( .A(n1311), .B(n1630), .Y(n1661) );
  AND2X1 U47 ( .A(n1630), .B(n1310), .Y(n1641) );
  AND2X1 U48 ( .A(n1311), .B(n1591), .Y(n1620) );
  AND2X1 U49 ( .A(n1591), .B(n1310), .Y(n1601) );
  AND2X1 U50 ( .A(n1311), .B(n940), .Y(n1581) );
  AND2X1 U51 ( .A(n940), .B(n1310), .Y(n1562) );
  OR2X1 U52 ( .A(n970), .B(n965), .Y(n968) );
  AND2X1 U53 ( .A(n1311), .B(n951), .Y(n1542) );
  OR2X1 U54 ( .A(n965), .B(n971), .Y(n966) );
  AND2X1 U55 ( .A(n1827), .B(\mem<32><0> ), .Y(n1491) );
  AND2X1 U56 ( .A(n1827), .B(\mem<32><1> ), .Y(n1503) );
  AND2X1 U57 ( .A(n1827), .B(\mem<32><2> ), .Y(n1336) );
  AND2X1 U58 ( .A(n1827), .B(\mem<32><3> ), .Y(n1349) );
  AND2X1 U59 ( .A(n1827), .B(\mem<32><4> ), .Y(n1362) );
  AND2X1 U60 ( .A(n1827), .B(\mem<32><5> ), .Y(n1375) );
  AND2X1 U61 ( .A(n1827), .B(\mem<32><6> ), .Y(n1388) );
  AND2X1 U62 ( .A(n1827), .B(\mem<32><7> ), .Y(n1401) );
  INVX1 U63 ( .A(rd1), .Y(n1014) );
  BUFX2 U64 ( .A(n961), .Y(n1010) );
  BUFX2 U65 ( .A(n961), .Y(n1009) );
  BUFX2 U66 ( .A(n960), .Y(n1007) );
  BUFX2 U67 ( .A(n960), .Y(n1006) );
  BUFX2 U68 ( .A(n959), .Y(n1004) );
  BUFX2 U69 ( .A(n959), .Y(n1003) );
  BUFX2 U70 ( .A(n958), .Y(n1001) );
  BUFX2 U71 ( .A(n958), .Y(n1000) );
  BUFX2 U72 ( .A(n957), .Y(n990) );
  BUFX2 U73 ( .A(n957), .Y(n989) );
  BUFX2 U74 ( .A(n956), .Y(n987) );
  BUFX2 U75 ( .A(n956), .Y(n986) );
  BUFX2 U76 ( .A(n955), .Y(n984) );
  BUFX2 U77 ( .A(n955), .Y(n983) );
  BUFX2 U78 ( .A(n954), .Y(n981) );
  BUFX2 U79 ( .A(n954), .Y(n980) );
  INVX1 U80 ( .A(\data_in_1c<0> ), .Y(n1028) );
  INVX1 U81 ( .A(\data_in_1c<1> ), .Y(n1029) );
  INVX1 U82 ( .A(\data_in_1c<2> ), .Y(n1030) );
  INVX1 U83 ( .A(\data_in_1c<3> ), .Y(n1031) );
  INVX1 U84 ( .A(\data_in_1c<4> ), .Y(n1032) );
  INVX1 U85 ( .A(\data_in_1c<5> ), .Y(n1033) );
  INVX1 U86 ( .A(\data_in_1c<6> ), .Y(n1034) );
  INVX1 U87 ( .A(\data_in_1c<7> ), .Y(n1035) );
  INVX1 U88 ( .A(\data_in_1c<8> ), .Y(n1036) );
  INVX1 U89 ( .A(\data_in_1c<9> ), .Y(n1037) );
  INVX1 U90 ( .A(\data_in_1c<10> ), .Y(n1038) );
  INVX1 U91 ( .A(\data_in_1c<11> ), .Y(n1039) );
  INVX1 U92 ( .A(\data_in_1c<12> ), .Y(n1040) );
  INVX1 U93 ( .A(\data_in_1c<13> ), .Y(n1041) );
  INVX1 U129 ( .A(\data_in_1c<14> ), .Y(n1042) );
  INVX1 U589 ( .A(\data_in_1c<15> ), .Y(n1043) );
  INVX1 U640 ( .A(wr), .Y(n1044) );
  INVX1 U659 ( .A(n1324), .Y(n1022) );
  INVX1 U660 ( .A(n1415), .Y(n1021) );
  INVX1 U664 ( .A(n1426), .Y(n1020) );
  INVX1 U666 ( .A(n1437), .Y(n1019) );
  INVX1 U672 ( .A(n1448), .Y(n1018) );
  INVX1 U675 ( .A(n1459), .Y(n1017) );
  INVX1 U679 ( .A(n1470), .Y(n1016) );
  INVX1 U682 ( .A(n1481), .Y(n1015) );
  AND2X1 U694 ( .A(wr1), .B(n1013), .Y(n1828) );
  INVX1 U697 ( .A(rst), .Y(n1013) );
  INVX2 U701 ( .A(n1013), .Y(n1012) );
  AND2X1 U706 ( .A(n387), .B(n372), .Y(n1) );
  INVX1 U712 ( .A(n1), .Y(n2) );
  AND2X1 U717 ( .A(n402), .B(n381), .Y(n3) );
  INVX1 U723 ( .A(n3), .Y(n4) );
  AND2X1 U728 ( .A(n1817), .B(n189), .Y(n5) );
  INVX1 U734 ( .A(n5), .Y(n6) );
  AND2X1 U739 ( .A(n973), .B(n289), .Y(n7) );
  INVX1 U745 ( .A(n7), .Y(n8) );
  OR2X1 U750 ( .A(n486), .B(n10), .Y(n9) );
  OR2X1 U756 ( .A(n473), .B(n474), .Y(n10) );
  OR2X1 U761 ( .A(n508), .B(n12), .Y(n11) );
  OR2X1 U767 ( .A(n487), .B(n507), .Y(n12) );
  OR2X1 U772 ( .A(n537), .B(n14), .Y(n13) );
  OR2X1 U786 ( .A(n522), .B(n523), .Y(n14) );
  OR2X1 U789 ( .A(n553), .B(n16), .Y(n15) );
  OR2X1 U801 ( .A(n538), .B(n552), .Y(n16) );
  OR2X1 U804 ( .A(n582), .B(n18), .Y(n17) );
  OR2X1 U816 ( .A(n567), .B(n568), .Y(n18) );
  OR2X1 U819 ( .A(n592), .B(n20), .Y(n19) );
  OR2X1 U831 ( .A(n583), .B(n591), .Y(n20) );
  OR2X1 U834 ( .A(n873), .B(n22), .Y(n21) );
  OR2X1 U846 ( .A(n871), .B(n872), .Y(n22) );
  OR2X1 U849 ( .A(n876), .B(n24), .Y(n23) );
  OR2X1 U861 ( .A(n874), .B(n875), .Y(n24) );
  OR2X1 U864 ( .A(n895), .B(n26), .Y(n25) );
  OR2X1 U870 ( .A(n893), .B(n894), .Y(n26) );
  OR2X1 U875 ( .A(n898), .B(n28), .Y(n27) );
  OR2X1 U882 ( .A(n896), .B(n897), .Y(n28) );
  OR2X1 U883 ( .A(n901), .B(n30), .Y(n29) );
  OR2X1 U884 ( .A(n899), .B(n900), .Y(n30) );
  OR2X1 U885 ( .A(n904), .B(n32), .Y(n31) );
  OR2X1 U886 ( .A(n902), .B(n903), .Y(n32) );
  OR2X1 U887 ( .A(n907), .B(n34), .Y(n33) );
  OR2X1 U888 ( .A(n905), .B(n906), .Y(n34) );
  OR2X1 U889 ( .A(n910), .B(n36), .Y(n35) );
  OR2X1 U890 ( .A(n908), .B(n909), .Y(n36) );
  OR2X1 U891 ( .A(n913), .B(n38), .Y(n37) );
  OR2X1 U892 ( .A(n911), .B(n912), .Y(n38) );
  OR2X1 U893 ( .A(n916), .B(n150), .Y(n50) );
  OR2X1 U894 ( .A(n914), .B(n915), .Y(n150) );
  AND2X1 U895 ( .A(n973), .B(n1828), .Y(n189) );
  AND2X1 U896 ( .A(n1828), .B(n1524), .Y(n289) );
  AND2X1 U897 ( .A(n940), .B(n942), .Y(n348) );
  INVX1 U898 ( .A(n348), .Y(n372) );
  AND2X1 U899 ( .A(n951), .B(n953), .Y(n379) );
  INVX1 U900 ( .A(n379), .Y(n381) );
  AND2X1 U901 ( .A(n940), .B(n941), .Y(n386) );
  INVX1 U902 ( .A(n386), .Y(n387) );
  AND2X1 U903 ( .A(n951), .B(n952), .Y(n401) );
  INVX1 U904 ( .A(n401), .Y(n402) );
  BUFX2 U905 ( .A(n1339), .Y(n408) );
  BUFX2 U906 ( .A(n1352), .Y(n409) );
  BUFX2 U907 ( .A(n1365), .Y(n421) );
  BUFX2 U908 ( .A(n1378), .Y(n422) );
  BUFX2 U909 ( .A(n1391), .Y(n434) );
  BUFX2 U910 ( .A(n1404), .Y(n435) );
  BUFX2 U911 ( .A(n1494), .Y(n447) );
  BUFX2 U912 ( .A(n1505), .Y(n448) );
  AND2X2 U913 ( .A(rd), .B(n1508), .Y(n460) );
  INVX1 U914 ( .A(n460), .Y(n461) );
  INVX1 U915 ( .A(n1314), .Y(n473) );
  INVX1 U916 ( .A(n1315), .Y(n474) );
  INVX1 U917 ( .A(n1316), .Y(n486) );
  INVX1 U918 ( .A(n1407), .Y(n487) );
  INVX1 U919 ( .A(n1408), .Y(n507) );
  INVX1 U920 ( .A(n1409), .Y(n508) );
  INVX1 U921 ( .A(n1418), .Y(n522) );
  INVX1 U922 ( .A(n1419), .Y(n523) );
  INVX1 U923 ( .A(n1420), .Y(n537) );
  INVX1 U924 ( .A(n1429), .Y(n538) );
  INVX1 U925 ( .A(n1430), .Y(n552) );
  INVX1 U926 ( .A(n1431), .Y(n553) );
  INVX1 U927 ( .A(n1440), .Y(n567) );
  INVX1 U928 ( .A(n1441), .Y(n568) );
  INVX1 U929 ( .A(n1442), .Y(n582) );
  INVX1 U930 ( .A(n1451), .Y(n583) );
  INVX1 U931 ( .A(n1452), .Y(n591) );
  INVX1 U932 ( .A(n1453), .Y(n592) );
  INVX1 U933 ( .A(n1462), .Y(n871) );
  INVX1 U934 ( .A(n1463), .Y(n872) );
  INVX1 U935 ( .A(n1464), .Y(n873) );
  INVX1 U936 ( .A(n1473), .Y(n874) );
  INVX1 U937 ( .A(n1474), .Y(n875) );
  INVX1 U938 ( .A(n1475), .Y(n876) );
  AND2X2 U939 ( .A(n1328), .B(n1327), .Y(n877) );
  INVX1 U940 ( .A(n877), .Y(n878) );
  AND2X2 U941 ( .A(n1341), .B(n1340), .Y(n879) );
  INVX1 U942 ( .A(n879), .Y(n880) );
  AND2X2 U943 ( .A(n1354), .B(n1353), .Y(n881) );
  INVX1 U944 ( .A(n881), .Y(n882) );
  AND2X2 U945 ( .A(n1367), .B(n1366), .Y(n883) );
  INVX1 U946 ( .A(n883), .Y(n884) );
  AND2X2 U947 ( .A(n1380), .B(n1379), .Y(n885) );
  INVX1 U948 ( .A(n885), .Y(n886) );
  AND2X2 U949 ( .A(n1393), .B(n1392), .Y(n887) );
  INVX1 U950 ( .A(n887), .Y(n888) );
  AND2X2 U951 ( .A(n1483), .B(n1482), .Y(n889) );
  INVX1 U952 ( .A(n889), .Y(n890) );
  AND2X2 U953 ( .A(n1496), .B(n1495), .Y(n891) );
  INVX1 U954 ( .A(n891), .Y(n892) );
  INVX1 U955 ( .A(n1321), .Y(n893) );
  INVX1 U956 ( .A(n1322), .Y(n894) );
  INVX1 U957 ( .A(n1323), .Y(n895) );
  INVX1 U958 ( .A(n1412), .Y(n896) );
  INVX1 U959 ( .A(n1413), .Y(n897) );
  INVX1 U960 ( .A(n1414), .Y(n898) );
  INVX1 U961 ( .A(n1423), .Y(n899) );
  INVX1 U962 ( .A(n1424), .Y(n900) );
  INVX1 U963 ( .A(n1425), .Y(n901) );
  INVX1 U964 ( .A(n1434), .Y(n902) );
  INVX1 U965 ( .A(n1435), .Y(n903) );
  INVX1 U966 ( .A(n1436), .Y(n904) );
  INVX1 U967 ( .A(n1445), .Y(n905) );
  INVX1 U968 ( .A(n1446), .Y(n906) );
  INVX1 U969 ( .A(n1447), .Y(n907) );
  INVX1 U970 ( .A(n1456), .Y(n908) );
  INVX1 U971 ( .A(n1457), .Y(n909) );
  INVX1 U972 ( .A(n1458), .Y(n910) );
  INVX1 U973 ( .A(n1467), .Y(n911) );
  INVX1 U974 ( .A(n1468), .Y(n912) );
  INVX1 U975 ( .A(n1469), .Y(n913) );
  INVX1 U976 ( .A(n1478), .Y(n914) );
  INVX1 U977 ( .A(n1479), .Y(n915) );
  INVX1 U978 ( .A(n1480), .Y(n916) );
  AND2X2 U979 ( .A(n1330), .B(n1329), .Y(n917) );
  INVX1 U980 ( .A(n917), .Y(n918) );
  AND2X2 U981 ( .A(n1343), .B(n1342), .Y(n919) );
  INVX1 U982 ( .A(n919), .Y(n920) );
  AND2X2 U983 ( .A(n1356), .B(n1355), .Y(n921) );
  INVX1 U984 ( .A(n921), .Y(n922) );
  AND2X2 U985 ( .A(n1369), .B(n1368), .Y(n923) );
  INVX1 U986 ( .A(n923), .Y(n924) );
  AND2X2 U987 ( .A(n1382), .B(n1381), .Y(n925) );
  INVX1 U988 ( .A(n925), .Y(n926) );
  AND2X2 U989 ( .A(n1395), .B(n1394), .Y(n927) );
  INVX1 U990 ( .A(n927), .Y(n928) );
  AND2X2 U991 ( .A(n1485), .B(n1484), .Y(n929) );
  INVX1 U992 ( .A(n929), .Y(n930) );
  AND2X2 U993 ( .A(n1498), .B(n1497), .Y(n931) );
  INVX1 U994 ( .A(n931), .Y(n932) );
  BUFX2 U995 ( .A(n1337), .Y(n933) );
  BUFX2 U996 ( .A(n1350), .Y(n934) );
  BUFX2 U997 ( .A(n1363), .Y(n935) );
  BUFX2 U998 ( .A(n1376), .Y(n936) );
  BUFX2 U999 ( .A(n1389), .Y(n937) );
  BUFX2 U1000 ( .A(n1402), .Y(n938) );
  BUFX2 U1001 ( .A(n1492), .Y(n939) );
  INVX1 U1002 ( .A(n970), .Y(n940) );
  INVX1 U1003 ( .A(n1499), .Y(n941) );
  INVX1 U1004 ( .A(n1500), .Y(n942) );
  BUFX2 U1005 ( .A(n1552), .Y(n970) );
  BUFX2 U1006 ( .A(n1838), .Y(err) );
  BUFX2 U1007 ( .A(n1335), .Y(n944) );
  BUFX2 U1008 ( .A(n1348), .Y(n945) );
  BUFX2 U1009 ( .A(n1361), .Y(n946) );
  BUFX2 U1010 ( .A(n1374), .Y(n947) );
  BUFX2 U1011 ( .A(n1387), .Y(n948) );
  BUFX2 U1012 ( .A(n1400), .Y(n949) );
  BUFX2 U1013 ( .A(n1490), .Y(n950) );
  INVX1 U1014 ( .A(n971), .Y(n951) );
  INVX1 U1015 ( .A(n1501), .Y(n952) );
  INVX1 U1016 ( .A(n1502), .Y(n953) );
  BUFX2 U1017 ( .A(n1514), .Y(n971) );
  BUFX2 U1018 ( .A(n1523), .Y(n972) );
  BUFX2 U1019 ( .A(n1541), .Y(n974) );
  BUFX2 U1020 ( .A(n1551), .Y(n975) );
  BUFX2 U1021 ( .A(n1561), .Y(n976) );
  BUFX2 U1022 ( .A(n1571), .Y(n977) );
  BUFX2 U1023 ( .A(n1580), .Y(n978) );
  BUFX2 U1024 ( .A(n1590), .Y(n979) );
  BUFX2 U1025 ( .A(n1610), .Y(n982) );
  BUFX2 U1026 ( .A(n1629), .Y(n985) );
  BUFX2 U1027 ( .A(n1650), .Y(n988) );
  BUFX2 U1028 ( .A(n1670), .Y(n991) );
  BUFX2 U1029 ( .A(n1679), .Y(n992) );
  BUFX2 U1030 ( .A(n1689), .Y(n993) );
  BUFX2 U1031 ( .A(n1698), .Y(n994) );
  BUFX2 U1032 ( .A(n1708), .Y(n995) );
  BUFX2 U1033 ( .A(n1717), .Y(n996) );
  BUFX2 U1034 ( .A(n1727), .Y(n997) );
  BUFX2 U1035 ( .A(n1736), .Y(n998) );
  BUFX2 U1036 ( .A(n1746), .Y(n999) );
  BUFX2 U1037 ( .A(n1765), .Y(n1002) );
  BUFX2 U1038 ( .A(n1785), .Y(n1005) );
  BUFX2 U1039 ( .A(n1805), .Y(n1008) );
  BUFX2 U1040 ( .A(n1818), .Y(n973) );
  AND2X1 U1041 ( .A(n1630), .B(n1318), .Y(n1817) );
  BUFX2 U1042 ( .A(n1837), .Y(n1011) );
  BUFX2 U1043 ( .A(n1600), .Y(n954) );
  BUFX2 U1044 ( .A(n1619), .Y(n955) );
  BUFX2 U1045 ( .A(n1640), .Y(n956) );
  BUFX2 U1046 ( .A(n1660), .Y(n957) );
  BUFX2 U1047 ( .A(n1755), .Y(n958) );
  BUFX2 U1048 ( .A(n1775), .Y(n959) );
  BUFX2 U1049 ( .A(n1795), .Y(n960) );
  BUFX2 U1050 ( .A(n1816), .Y(n961) );
  AND2X1 U1051 ( .A(enable), .B(n1013), .Y(n962) );
  INVX1 U1052 ( .A(n962), .Y(n963) );
  AND2X1 U1053 ( .A(n1513), .B(n1512), .Y(n964) );
  INVX1 U1054 ( .A(n964), .Y(n965) );
  INVX1 U1055 ( .A(n966), .Y(n967) );
  INVX1 U1056 ( .A(n968), .Y(n969) );
  AND2X1 U1057 ( .A(n951), .B(n1310), .Y(n1524) );
endmodule


module dff_216 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_217 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_218 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_219 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_212 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_213 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_214 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_215 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_208 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_209 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_210 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_211 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module mem_state_reg ( clk, rst, .state({\state<3> , \state<2> , \state<1> , 
        \state<0> }), .next_state({\next_state<3> , \next_state<2> , 
        \next_state<1> , \next_state<0> }) );
  input clk, rst, \state<3> , \state<2> , \state<1> , \state<0> ;
  output \next_state<3> , \next_state<2> , \next_state<1> , \next_state<0> ;


  dff_0 \STATE[0]  ( .q(), .d(\next_state<0> ), .clk(clk), .rst(rst) );
  dff_1 \STATE[1]  ( .q(), .d(\next_state<1> ), .clk(clk), .rst(rst) );
  dff_2 \STATE[2]  ( .q(), .d(\next_state<2> ), .clk(clk), .rst(rst) );
  dff_3 \STATE[3]  ( .q(), .d(\next_state<3> ), .clk(clk), .rst(rst) );
endmodule


module mem_next_state ( rd, wr, hit, dirty, .state({\state<3> , \state<2> , 
        \state<1> , \state<0> }), err, .next_state({\next_state<3> , 
        \next_state<2> , \next_state<1> , \next_state<0> }) );
  input rd, wr, hit, dirty, \state<3> , \state<2> , \state<1> , \state<0> ;
  output err, \next_state<3> , \next_state<2> , \next_state<1> ,
         \next_state<0> ;
  wire   n18, n19, n20, n21, n22, n23, n24, n25, n26, n29, n32, n33, n34, n35,
         n36, n37, n39, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n27, n28, n30, n31, n38, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52;

  NAND3X1 U21 ( .A(n12), .B(n27), .C(n8), .Y(\next_state<3> ) );
  AOI21X1 U22 ( .A(n31), .B(n19), .C(n20), .Y(n18) );
  NAND3X1 U23 ( .A(n3), .B(n13), .C(n7), .Y(\next_state<2> ) );
  AOI21X1 U24 ( .A(n16), .B(n25), .C(n26), .Y(n23) );
  OAI21X1 U25 ( .A(n30), .B(n38), .C(n12), .Y(n26) );
  AOI22X1 U27 ( .A(n16), .B(n42), .C(n29), .D(n19), .Y(n21) );
  AOI21X1 U28 ( .A(n52), .B(n51), .C(dirty), .Y(n24) );
  NAND3X1 U29 ( .A(n30), .B(n41), .C(n47), .Y(\next_state<1> ) );
  OAI21X1 U30 ( .A(n15), .B(n30), .C(n1), .Y(n20) );
  AOI21X1 U31 ( .A(n40), .B(n14), .C(err), .Y(n32) );
  NAND3X1 U33 ( .A(n2), .B(n6), .C(n44), .Y(\next_state<0> ) );
  NAND3X1 U34 ( .A(n13), .B(n27), .C(n41), .Y(n35) );
  AOI21X1 U37 ( .A(n9), .B(n31), .C(n36), .Y(n22) );
  OAI21X1 U38 ( .A(n38), .B(n41), .C(n46), .Y(n36) );
  AOI22X1 U41 ( .A(rd), .B(n42), .C(wr), .D(n42), .Y(n34) );
  NAND3X1 U42 ( .A(n9), .B(n43), .C(n29), .Y(n37) );
  AOI22X1 U43 ( .A(rd), .B(n25), .C(wr), .D(n25), .Y(n33) );
  AND2X1 U1 ( .A(\state<2> ), .B(\state<3> ), .Y(n39) );
  INVX1 U2 ( .A(hit), .Y(n43) );
  INVX1 U3 ( .A(wr), .Y(n52) );
  INVX1 U4 ( .A(\state<3> ), .Y(n45) );
  INVX1 U5 ( .A(\state<2> ), .Y(n48) );
  INVX1 U6 ( .A(\state<0> ), .Y(n50) );
  INVX1 U7 ( .A(\state<1> ), .Y(n49) );
  AND2X1 U8 ( .A(n39), .B(n43), .Y(n25) );
  AND2X1 U9 ( .A(n39), .B(n10), .Y(err) );
  AND2X1 U10 ( .A(n45), .B(n48), .Y(n29) );
  INVX1 U11 ( .A(rd), .Y(n51) );
  AND2X1 U12 ( .A(\state<1> ), .B(\state<0> ), .Y(n19) );
  INVX1 U13 ( .A(n20), .Y(n47) );
  INVX1 U14 ( .A(err), .Y(n46) );
  BUFX2 U15 ( .A(n32), .Y(n1) );
  BUFX2 U16 ( .A(n33), .Y(n2) );
  BUFX2 U17 ( .A(n21), .Y(n3) );
  BUFX2 U18 ( .A(n37), .Y(n4) );
  INVX1 U19 ( .A(n4), .Y(n42) );
  BUFX2 U20 ( .A(n35), .Y(n5) );
  INVX1 U26 ( .A(n5), .Y(n44) );
  BUFX2 U32 ( .A(n34), .Y(n6) );
  BUFX2 U35 ( .A(n23), .Y(n7) );
  BUFX2 U36 ( .A(n18), .Y(n8) );
  AND2X1 U39 ( .A(n49), .B(n50), .Y(n9) );
  INVX1 U40 ( .A(n9), .Y(n10) );
  AND2X1 U44 ( .A(\state<3> ), .B(n19), .Y(n11) );
  INVX1 U45 ( .A(n11), .Y(n12) );
  BUFX2 U46 ( .A(n22), .Y(n13) );
  AND2X1 U47 ( .A(\state<3> ), .B(n48), .Y(n14) );
  INVX1 U48 ( .A(n14), .Y(n15) );
  BUFX2 U49 ( .A(n24), .Y(n16) );
  AND2X1 U50 ( .A(n9), .B(n14), .Y(n17) );
  INVX1 U51 ( .A(n17), .Y(n27) );
  AND2X1 U52 ( .A(\state<0> ), .B(n49), .Y(n28) );
  INVX1 U53 ( .A(n28), .Y(n30) );
  AND2X1 U54 ( .A(\state<2> ), .B(n45), .Y(n31) );
  INVX1 U55 ( .A(n31), .Y(n38) );
  AND2X1 U56 ( .A(\state<1> ), .B(n50), .Y(n40) );
  INVX1 U57 ( .A(n40), .Y(n41) );
endmodule


module mem_signals ( hit, .state({\state<3> , \state<2> , \state<1> , 
        \state<0> }), stall, done, cache_wr, cache_hit, .cache_offset({
        \cache_offset<1> , \cache_offset<0> }), cache_sel, comp, mem_wr, 
        mem_rd, .mem_offset({\mem_offset<1> , \mem_offset<0> }), mem_sel );
  input hit, \state<3> , \state<2> , \state<1> , \state<0> ;
  output stall, done, cache_wr, cache_hit, \cache_offset<1> ,
         \cache_offset<0> , cache_sel, comp, mem_wr, mem_rd, \mem_offset<1> ,
         \mem_offset<0> , mem_sel;
  wire   n51, n13, n18, n19, n20, n23, n26, n27, n28, n29, n30, n32, n34, n1,
         n2, n3, n4, n5, n6, n8, n9, n10, n11, n12, n14, n15, n16, n17, n21,
         n22, n24, n25, n31, n33, n35, n36, n37, n38, n39, n40, n41, n42, n46,
         n47, n48, n49, n50;

  NAND3X1 U17 ( .A(n13), .B(n40), .C(n31), .Y(stall) );
  OAI21X1 U18 ( .A(n35), .B(n21), .C(n2), .Y(mem_wr) );
  NAND3X1 U19 ( .A(n47), .B(n46), .C(n25), .Y(n18) );
  OAI21X1 U20 ( .A(n19), .B(n40), .C(n15), .Y(mem_sel) );
  OAI21X1 U21 ( .A(n19), .B(n40), .C(n6), .Y(\mem_offset<1> ) );
  XNOR2X1 U23 ( .A(n14), .B(n46), .Y(n23) );
  OAI21X1 U25 ( .A(n35), .B(n24), .C(n16), .Y(done) );
  AOI22X1 U26 ( .A(n22), .B(n28), .C(n17), .D(n37), .Y(n27) );
  NAND3X1 U27 ( .A(n15), .B(n40), .C(n9), .Y(n51) );
  AOI22X1 U28 ( .A(n22), .B(n30), .C(n37), .D(n48), .Y(n29) );
  NAND3X1 U30 ( .A(n25), .B(n46), .C(\state<2> ), .Y(n20) );
  OAI21X1 U32 ( .A(n48), .B(n36), .C(n1), .Y(cache_sel) );
  AOI21X1 U33 ( .A(n17), .B(n36), .C(n41), .Y(n32) );
  OAI21X1 U34 ( .A(n48), .B(n40), .C(n4), .Y(\cache_offset<1> ) );
  OAI21X1 U36 ( .A(\state<2> ), .B(n39), .C(n35), .Y(n28) );
  XNOR2X1 U39 ( .A(n11), .B(n47), .Y(n34) );
  NAND3X1 U41 ( .A(n17), .B(n37), .C(hit), .Y(n26) );
  XNOR2X1 U45 ( .A(\state<0> ), .B(n49), .Y(n19) );
  OR2X1 U1 ( .A(n39), .B(n47), .Y(n30) );
  AND2X1 U2 ( .A(n34), .B(n50), .Y(\cache_offset<0> ) );
  INVX1 U3 ( .A(n19), .Y(n48) );
  INVX1 U4 ( .A(\state<0> ), .Y(n50) );
  INVX1 U5 ( .A(\state<1> ), .Y(n49) );
  INVX1 U6 ( .A(\state<3> ), .Y(n46) );
  INVX1 U7 ( .A(\state<2> ), .Y(n47) );
  AND2X1 U8 ( .A(n23), .B(n50), .Y(\mem_offset<0> ) );
  OR2X1 U9 ( .A(n35), .B(\state<3> ), .Y(n13) );
  BUFX2 U10 ( .A(n32), .Y(n1) );
  BUFX2 U11 ( .A(n18), .Y(n2) );
  AND2X1 U12 ( .A(n17), .B(n28), .Y(n3) );
  INVX1 U13 ( .A(n3), .Y(n4) );
  AND2X1 U14 ( .A(n17), .B(n36), .Y(n5) );
  INVX1 U15 ( .A(n5), .Y(n6) );
  BUFX2 U16 ( .A(n51), .Y(cache_wr) );
  BUFX2 U22 ( .A(n27), .Y(n8) );
  INVX1 U24 ( .A(n8), .Y(comp) );
  BUFX2 U29 ( .A(n29), .Y(n9) );
  AND2X1 U31 ( .A(n46), .B(n49), .Y(n10) );
  INVX1 U35 ( .A(n10), .Y(n11) );
  AND2X1 U37 ( .A(n47), .B(n49), .Y(n12) );
  INVX1 U38 ( .A(n12), .Y(n14) );
  BUFX2 U40 ( .A(n20), .Y(n15) );
  INVX1 U42 ( .A(cache_hit), .Y(n16) );
  INVX1 U43 ( .A(n26), .Y(cache_hit) );
  AND2X1 U44 ( .A(n48), .B(n46), .Y(n17) );
  INVX1 U46 ( .A(n17), .Y(n21) );
  AND2X1 U47 ( .A(\state<3> ), .B(n48), .Y(n22) );
  INVX1 U48 ( .A(n22), .Y(n24) );
  INVX1 U49 ( .A(n31), .Y(n25) );
  AND2X1 U50 ( .A(n48), .B(n39), .Y(n31) );
  AND2X1 U51 ( .A(\state<2> ), .B(n39), .Y(n33) );
  INVX1 U52 ( .A(n33), .Y(n35) );
  INVX1 U53 ( .A(n37), .Y(n36) );
  AND2X1 U54 ( .A(n47), .B(n39), .Y(n37) );
  AND2X1 U55 ( .A(\state<1> ), .B(\state<0> ), .Y(n38) );
  INVX1 U56 ( .A(n38), .Y(n39) );
  INVX1 U57 ( .A(n41), .Y(n40) );
  AND2X1 U58 ( .A(\state<3> ), .B(n37), .Y(n41) );
  INVX1 U59 ( .A(n42), .Y(mem_rd) );
  INVX1 U60 ( .A(mem_sel), .Y(n42) );
endmodule


module cache_cache_id0 ( enable, clk, rst, createdump, .tag_in({\tag_in<4> , 
        \tag_in<3> , \tag_in<2> , \tag_in<1> , \tag_in<0> }), .index({
        \index<7> , \index<6> , \index<5> , \index<4> , \index<3> , \index<2> , 
        \index<1> , \index<0> }), .offset({\offset<2> , \offset<1> , 
        \offset<0> }), .data_in({\data_in<15> , \data_in<14> , \data_in<13> , 
        \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> , 
        \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , 
        \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), comp, write, 
        valid_in, .tag_out({\tag_out<4> , \tag_out<3> , \tag_out<2> , 
        \tag_out<1> , \tag_out<0> }), .data_out({\data_out<15> , 
        \data_out<14> , \data_out<13> , \data_out<12> , \data_out<11> , 
        \data_out<10> , \data_out<9> , \data_out<8> , \data_out<7> , 
        \data_out<6> , \data_out<5> , \data_out<4> , \data_out<3> , 
        \data_out<2> , \data_out<1> , \data_out<0> }), hit, dirty, valid, err
 );
  input enable, clk, rst, createdump, \tag_in<4> , \tag_in<3> , \tag_in<2> ,
         \tag_in<1> , \tag_in<0> , \index<7> , \index<6> , \index<5> ,
         \index<4> , \index<3> , \index<2> , \index<1> , \index<0> ,
         \offset<2> , \offset<1> , \offset<0> , \data_in<15> , \data_in<14> ,
         \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> ,
         \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> ,
         \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> ,
         comp, write, valid_in;
  output \tag_out<4> , \tag_out<3> , \tag_out<2> , \tag_out<1> , \tag_out<0> ,
         \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , hit,
         dirty, valid, err;
  wire   n188, n189, n190, n191, \w0<15> , \w0<14> , \w0<13> , \w0<12> ,
         \w0<11> , \w0<10> , \w0<9> , \w0<8> , \w0<7> , \w0<6> , \w0<5> ,
         \w0<4> , \w0<3> , \w0<2> , \w0<1> , \w0<0> , \w1<15> , \w1<14> ,
         \w1<13> , \w1<12> , \w1<11> , \w1<10> , \w1<9> , \w1<8> , \w1<7> ,
         \w1<6> , \w1<5> , \w1<4> , \w1<3> , \w1<2> , \w1<1> , \w1<0> ,
         \w2<15> , \w2<14> , \w2<13> , \w2<12> , \w2<11> , \w2<10> , \w2<9> ,
         \w2<8> , \w2<7> , \w2<6> , \w2<5> , \w2<4> , \w2<3> , \w2<2> ,
         \w2<1> , \w2<0> , \w3<15> , \w3<14> , \w3<13> , \w3<12> , \w3<11> ,
         \w3<10> , \w3<9> , \w3<8> , \w3<7> , \w3<6> , \w3<5> , \w3<4> ,
         \w3<3> , \w3<2> , \w3<1> , \w3<0> , dirtybit, validbit, n17, n1, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n15, n18, n20, n22, n24,
         n26, n28, n30, n32, n34, n36, n38, n40, n42, n44, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n187;

  NAND3X1 U21 ( .A(n104), .B(n50), .C(validbit), .Y(n17) );
  memc_Size16_3 mem_w0 ( .data_out({\w0<15> , \w0<14> , \w0<13> , \w0<12> , 
        \w0<11> , \w0<10> , \w0<9> , \w0<8> , \w0<7> , \w0<6> , \w0<5> , 
        \w0<4> , \w0<3> , \w0<2> , \w0<1> , \w0<0> }), .addr({\index<7> , 
        \index<6> , \index<5> , n137, n135, n133, n131, n1}), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), .write(n12), .clk(clk), .rst(n129), 
        .createdump(createdump), .file_id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  memc_Size16_2 mem_w1 ( .data_out({\w1<15> , \w1<14> , \w1<13> , \w1<12> , 
        \w1<11> , \w1<10> , \w1<9> , \w1<8> , \w1<7> , \w1<6> , \w1<5> , 
        \w1<4> , \w1<3> , \w1<2> , \w1<1> , \w1<0> }), .addr({\index<7> , 
        \index<6> , \index<5> , n137, n135, n133, n131, n1}), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), .write(n10), .clk(clk), .rst(n129), 
        .createdump(createdump), .file_id({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}) );
  memc_Size16_1 mem_w2 ( .data_out({\w2<15> , \w2<14> , \w2<13> , \w2<12> , 
        \w2<11> , \w2<10> , \w2<9> , \w2<8> , \w2<7> , \w2<6> , \w2<5> , 
        \w2<4> , \w2<3> , \w2<2> , \w2<1> , \w2<0> }), .addr({\index<7> , 
        \index<6> , \index<5> , n137, n135, n133, n131, n1}), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), .write(n8), .clk(clk), .rst(n129), 
        .createdump(createdump), .file_id({1'b0, 1'b0, 1'b0, 1'b1, 1'b0}) );
  memc_Size16_0 mem_w3 ( .data_out({\w3<15> , \w3<14> , \w3<13> , \w3<12> , 
        \w3<11> , \w3<10> , \w3<9> , \w3<8> , \w3<7> , \w3<6> , \w3<5> , 
        \w3<4> , \w3<3> , \w3<2> , \w3<1> , \w3<0> }), .addr({\index<7> , 
        \index<6> , \index<5> , n137, n135, n133, n131, n1}), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), .write(n6), .clk(clk), .rst(n129), 
        .createdump(createdump), .file_id({1'b0, 1'b0, 1'b0, 1'b1, 1'b1}) );
  memc_Size5 mem_tg ( .data_out({\tag_out<4> , n188, n189, n190, n191}), 
        .addr({\index<7> , \index<6> , \index<5> , n137, n135, n133, n131, 
        \index<0> }), .data_in({\tag_in<4> , \tag_in<3> , \tag_in<2> , 
        \tag_in<1> , \tag_in<0> }), .write(n114), .clk(clk), .rst(n129), 
        .createdump(createdump), .file_id({1'b0, 1'b0, 1'b1, 1'b0, 1'b0}) );
  memc_Size1 mem_dr ( .data_out(dirtybit), .addr({\index<7> , \index<6> , 
        \index<5> , n137, n135, n133, n131, n1}), .data_in(comp), .write(n128), 
        .clk(clk), .rst(n129), .createdump(createdump), .file_id({1'b0, 1'b0, 
        1'b1, 1'b0, 1'b1}) );
  memv mem_vl ( .data_out(validbit), .addr({\index<7> , \index<6> , \index<5> , 
        n137, n135, n133, n131, n1}), .data_in(valid_in), .write(n113), .clk(
        clk), .rst(n129), .createdump(createdump), .file_id({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}) );
  INVX1 U3 ( .A(\tag_in<1> ), .Y(n125) );
  INVX1 U4 ( .A(\tag_in<3> ), .Y(n126) );
  INVX1 U5 ( .A(\index<4> ), .Y(n138) );
  INVX1 U6 ( .A(\tag_in<0> ), .Y(n123) );
  INVX1 U7 ( .A(\tag_in<2> ), .Y(n127) );
  INVX1 U8 ( .A(comp), .Y(n139) );
  INVX1 U9 ( .A(\offset<1> ), .Y(n148) );
  INVX1 U10 ( .A(\index<2> ), .Y(n134) );
  BUFX2 U11 ( .A(\index<0> ), .Y(n1) );
  BUFX2 U12 ( .A(n188), .Y(\tag_out<3> ) );
  INVX4 U13 ( .A(n132), .Y(n131) );
  AND2X2 U14 ( .A(enable), .B(n130), .Y(n104) );
  INVX1 U15 ( .A(n146), .Y(n3) );
  AND2X1 U16 ( .A(write), .B(n139), .Y(n49) );
  INVX1 U17 ( .A(write), .Y(n146) );
  INVX1 U18 ( .A(n46), .Y(n4) );
  INVX1 U19 ( .A(\index<1> ), .Y(n132) );
  AND2X2 U20 ( .A(n49), .B(n104), .Y(n114) );
  OR2X2 U22 ( .A(n145), .B(n112), .Y(n5) );
  INVX1 U23 ( .A(n5), .Y(n6) );
  OR2X2 U24 ( .A(n145), .B(n98), .Y(n7) );
  INVX1 U25 ( .A(n7), .Y(n8) );
  OR2X2 U26 ( .A(n145), .B(n100), .Y(n9) );
  INVX1 U27 ( .A(n9), .Y(n10) );
  OR2X2 U28 ( .A(n145), .B(n105), .Y(n11) );
  INVX1 U29 ( .A(n11), .Y(n12) );
  AND2X2 U30 ( .A(n71), .B(n53), .Y(n13) );
  INVX1 U31 ( .A(n13), .Y(\data_out<0> ) );
  AND2X2 U32 ( .A(n72), .B(n54), .Y(n15) );
  INVX1 U33 ( .A(n15), .Y(\data_out<1> ) );
  AND2X2 U34 ( .A(n55), .B(n73), .Y(n18) );
  INVX1 U35 ( .A(n18), .Y(\data_out<2> ) );
  AND2X2 U36 ( .A(n74), .B(n56), .Y(n20) );
  INVX1 U37 ( .A(n20), .Y(\data_out<3> ) );
  AND2X2 U38 ( .A(n75), .B(n57), .Y(n22) );
  INVX1 U39 ( .A(n22), .Y(\data_out<4> ) );
  AND2X2 U40 ( .A(n76), .B(n58), .Y(n24) );
  INVX1 U41 ( .A(n24), .Y(\data_out<5> ) );
  AND2X2 U42 ( .A(n77), .B(n59), .Y(n26) );
  INVX1 U43 ( .A(n26), .Y(\data_out<6> ) );
  AND2X2 U44 ( .A(n78), .B(n60), .Y(n28) );
  INVX1 U45 ( .A(n28), .Y(\data_out<7> ) );
  AND2X2 U46 ( .A(n79), .B(n61), .Y(n30) );
  INVX1 U47 ( .A(n30), .Y(\data_out<8> ) );
  AND2X2 U48 ( .A(n80), .B(n62), .Y(n32) );
  INVX1 U49 ( .A(n32), .Y(\data_out<9> ) );
  AND2X2 U50 ( .A(n81), .B(n63), .Y(n34) );
  INVX1 U51 ( .A(n34), .Y(\data_out<10> ) );
  AND2X2 U52 ( .A(n82), .B(n64), .Y(n36) );
  INVX1 U53 ( .A(n36), .Y(\data_out<11> ) );
  AND2X2 U54 ( .A(n83), .B(n65), .Y(n38) );
  INVX1 U55 ( .A(n38), .Y(\data_out<12> ) );
  AND2X2 U56 ( .A(n84), .B(n66), .Y(n40) );
  INVX1 U57 ( .A(n40), .Y(\data_out<13> ) );
  AND2X2 U58 ( .A(n85), .B(n67), .Y(n42) );
  INVX1 U59 ( .A(n42), .Y(\data_out<14> ) );
  AND2X2 U60 ( .A(n86), .B(n68), .Y(n44) );
  INVX1 U61 ( .A(n44), .Y(\data_out<15> ) );
  OR2X2 U62 ( .A(n48), .B(n47), .Y(n46) );
  OR2X2 U63 ( .A(n51), .B(n52), .Y(n47) );
  AND2X2 U64 ( .A(n88), .B(n70), .Y(n48) );
  INVX1 U65 ( .A(n49), .Y(n50) );
  OR2X2 U66 ( .A(n141), .B(n140), .Y(n51) );
  OR2X2 U67 ( .A(n143), .B(n142), .Y(n52) );
  BUFX2 U68 ( .A(n151), .Y(n53) );
  BUFX2 U69 ( .A(n153), .Y(n54) );
  BUFX2 U70 ( .A(n155), .Y(n55) );
  BUFX2 U71 ( .A(n157), .Y(n56) );
  BUFX2 U72 ( .A(n159), .Y(n57) );
  BUFX2 U73 ( .A(n161), .Y(n58) );
  BUFX2 U74 ( .A(n163), .Y(n59) );
  BUFX2 U75 ( .A(n165), .Y(n60) );
  BUFX2 U76 ( .A(n167), .Y(n61) );
  BUFX2 U77 ( .A(n169), .Y(n62) );
  BUFX2 U78 ( .A(n171), .Y(n63) );
  BUFX2 U79 ( .A(n173), .Y(n64) );
  BUFX2 U80 ( .A(n175), .Y(n65) );
  BUFX2 U81 ( .A(n177), .Y(n66) );
  BUFX2 U82 ( .A(n179), .Y(n67) );
  BUFX2 U83 ( .A(n183), .Y(n68) );
  AND2X2 U84 ( .A(n120), .B(n121), .Y(n69) );
  INVX1 U85 ( .A(n69), .Y(n70) );
  BUFX2 U86 ( .A(n152), .Y(n71) );
  BUFX2 U87 ( .A(n154), .Y(n72) );
  BUFX2 U88 ( .A(n156), .Y(n73) );
  BUFX2 U89 ( .A(n158), .Y(n74) );
  BUFX2 U90 ( .A(n160), .Y(n75) );
  BUFX2 U91 ( .A(n162), .Y(n76) );
  BUFX2 U92 ( .A(n164), .Y(n77) );
  BUFX2 U93 ( .A(n166), .Y(n78) );
  BUFX2 U94 ( .A(n168), .Y(n79) );
  BUFX2 U95 ( .A(n170), .Y(n80) );
  BUFX2 U96 ( .A(n172), .Y(n81) );
  BUFX2 U97 ( .A(n174), .Y(n82) );
  BUFX2 U98 ( .A(n176), .Y(n83) );
  BUFX2 U99 ( .A(n178), .Y(n84) );
  BUFX2 U100 ( .A(n180), .Y(n85) );
  BUFX2 U101 ( .A(n184), .Y(n86) );
  AND2X2 U102 ( .A(\tag_in<4> ), .B(\tag_out<4> ), .Y(n87) );
  INVX1 U103 ( .A(n87), .Y(n88) );
  AND2X2 U104 ( .A(n104), .B(n4), .Y(n89) );
  INVX1 U105 ( .A(n89), .Y(n90) );
  AND2X2 U106 ( .A(n104), .B(n144), .Y(n91) );
  INVX1 U107 ( .A(n91), .Y(n92) );
  INVX1 U108 ( .A(n91), .Y(n93) );
  AND2X1 U109 ( .A(n150), .B(n95), .Y(n94) );
  AND2X1 U110 ( .A(\offset<1> ), .B(n96), .Y(n95) );
  AND2X1 U111 ( .A(n146), .B(n104), .Y(n96) );
  AND2X1 U112 ( .A(\offset<2> ), .B(n148), .Y(n97) );
  INVX1 U113 ( .A(n97), .Y(n98) );
  AND2X1 U114 ( .A(n150), .B(\offset<1> ), .Y(n99) );
  INVX1 U115 ( .A(n99), .Y(n100) );
  BUFX2 U116 ( .A(n187), .Y(dirty) );
  AND2X2 U117 ( .A(dirtybit), .B(n104), .Y(n102) );
  INVX1 U118 ( .A(n102), .Y(n103) );
  INVX1 U119 ( .A(n17), .Y(valid) );
  OR2X1 U120 ( .A(\offset<1> ), .B(\offset<2> ), .Y(n105) );
  AND2X1 U121 ( .A(comp), .B(n124), .Y(n106) );
  INVX1 U122 ( .A(n106), .Y(n107) );
  BUFX2 U123 ( .A(n147), .Y(n108) );
  INVX1 U124 ( .A(n108), .Y(n181) );
  BUFX2 U125 ( .A(n149), .Y(n109) );
  INVX1 U126 ( .A(n109), .Y(n182) );
  INVX1 U127 ( .A(\offset<2> ), .Y(n150) );
  AND2X1 U128 ( .A(n111), .B(n96), .Y(n110) );
  AND2X1 U129 ( .A(\offset<2> ), .B(\offset<1> ), .Y(n111) );
  INVX1 U130 ( .A(n111), .Y(n112) );
  INVX1 U131 ( .A(n115), .Y(n113) );
  INVX1 U132 ( .A(n114), .Y(n115) );
  INVX1 U133 ( .A(n116), .Y(err) );
  INVX1 U134 ( .A(\offset<0> ), .Y(n116) );
  BUFX2 U135 ( .A(n191), .Y(\tag_out<0> ) );
  BUFX2 U136 ( .A(n190), .Y(\tag_out<1> ) );
  INVX1 U137 ( .A(\tag_in<4> ), .Y(n120) );
  INVX1 U138 ( .A(\tag_out<4> ), .Y(n121) );
  BUFX2 U139 ( .A(n189), .Y(\tag_out<2> ) );
  XNOR2X1 U140 ( .A(n191), .B(n123), .Y(n142) );
  BUFX2 U141 ( .A(n46), .Y(n124) );
  XNOR2X1 U142 ( .A(n190), .B(n125), .Y(n143) );
  XNOR2X1 U143 ( .A(n188), .B(n126), .Y(n140) );
  XNOR2X1 U144 ( .A(n189), .B(n127), .Y(n141) );
  OAI21X1 U145 ( .A(n92), .B(n146), .C(n115), .Y(n128) );
  INVX1 U146 ( .A(n93), .Y(hit) );
  INVX1 U147 ( .A(n46), .Y(n144) );
  INVX8 U148 ( .A(n130), .Y(n129) );
  INVX8 U149 ( .A(rst), .Y(n130) );
  INVX8 U150 ( .A(n134), .Y(n133) );
  INVX8 U151 ( .A(n136), .Y(n135) );
  INVX8 U152 ( .A(\index<3> ), .Y(n136) );
  INVX8 U153 ( .A(n138), .Y(n137) );
  OAI21X1 U154 ( .A(n146), .B(n90), .C(n115), .Y(n185) );
  INVX2 U155 ( .A(n185), .Y(n145) );
  AOI21X1 U156 ( .A(n3), .B(n107), .C(n103), .Y(n187) );
  NAND3X1 U157 ( .A(\offset<2> ), .B(n96), .C(n148), .Y(n147) );
  AOI22X1 U158 ( .A(n181), .B(\w2<0> ), .C(n110), .D(\w3<0> ), .Y(n152) );
  NAND3X1 U159 ( .A(n148), .B(n96), .C(n150), .Y(n149) );
  AOI22X1 U160 ( .A(n182), .B(\w0<0> ), .C(\w1<0> ), .D(n94), .Y(n151) );
  AOI22X1 U161 ( .A(n181), .B(\w2<1> ), .C(\w3<1> ), .D(n110), .Y(n154) );
  AOI22X1 U162 ( .A(n182), .B(\w0<1> ), .C(\w1<1> ), .D(n94), .Y(n153) );
  AOI22X1 U163 ( .A(n181), .B(\w2<2> ), .C(n110), .D(\w3<2> ), .Y(n156) );
  AOI22X1 U164 ( .A(n182), .B(\w0<2> ), .C(n94), .D(\w1<2> ), .Y(n155) );
  AOI22X1 U165 ( .A(n181), .B(\w2<3> ), .C(\w3<3> ), .D(n110), .Y(n158) );
  AOI22X1 U166 ( .A(n182), .B(\w0<3> ), .C(\w1<3> ), .D(n94), .Y(n157) );
  AOI22X1 U167 ( .A(n181), .B(\w2<4> ), .C(\w3<4> ), .D(n110), .Y(n160) );
  AOI22X1 U168 ( .A(n182), .B(\w0<4> ), .C(\w1<4> ), .D(n94), .Y(n159) );
  AOI22X1 U169 ( .A(n181), .B(\w2<5> ), .C(\w3<5> ), .D(n110), .Y(n162) );
  AOI22X1 U170 ( .A(n182), .B(\w0<5> ), .C(\w1<5> ), .D(n94), .Y(n161) );
  AOI22X1 U171 ( .A(n181), .B(\w2<6> ), .C(\w3<6> ), .D(n110), .Y(n164) );
  AOI22X1 U172 ( .A(n182), .B(\w0<6> ), .C(\w1<6> ), .D(n94), .Y(n163) );
  AOI22X1 U173 ( .A(n181), .B(\w2<7> ), .C(n110), .D(\w3<7> ), .Y(n166) );
  AOI22X1 U174 ( .A(n182), .B(\w0<7> ), .C(\w1<7> ), .D(n94), .Y(n165) );
  AOI22X1 U175 ( .A(n181), .B(\w2<8> ), .C(n110), .D(\w3<8> ), .Y(n168) );
  AOI22X1 U176 ( .A(n182), .B(\w0<8> ), .C(\w1<8> ), .D(n94), .Y(n167) );
  AOI22X1 U177 ( .A(n181), .B(\w2<9> ), .C(\w3<9> ), .D(n110), .Y(n170) );
  AOI22X1 U178 ( .A(n182), .B(\w0<9> ), .C(n94), .D(\w1<9> ), .Y(n169) );
  AOI22X1 U179 ( .A(n181), .B(\w2<10> ), .C(n110), .D(\w3<10> ), .Y(n172) );
  AOI22X1 U180 ( .A(n182), .B(\w0<10> ), .C(\w1<10> ), .D(n94), .Y(n171) );
  AOI22X1 U181 ( .A(n181), .B(\w2<11> ), .C(n110), .D(\w3<11> ), .Y(n174) );
  AOI22X1 U182 ( .A(n182), .B(\w0<11> ), .C(\w1<11> ), .D(n94), .Y(n173) );
  AOI22X1 U183 ( .A(n181), .B(\w2<12> ), .C(n110), .D(\w3<12> ), .Y(n176) );
  AOI22X1 U184 ( .A(n182), .B(\w0<12> ), .C(\w1<12> ), .D(n94), .Y(n175) );
  AOI22X1 U185 ( .A(n181), .B(\w2<13> ), .C(\w3<13> ), .D(n110), .Y(n178) );
  AOI22X1 U186 ( .A(n182), .B(\w0<13> ), .C(\w1<13> ), .D(n94), .Y(n177) );
  AOI22X1 U187 ( .A(n181), .B(\w2<14> ), .C(n110), .D(\w3<14> ), .Y(n180) );
  AOI22X1 U188 ( .A(n182), .B(\w0<14> ), .C(n94), .D(\w1<14> ), .Y(n179) );
  AOI22X1 U189 ( .A(n181), .B(\w2<15> ), .C(n110), .D(\w3<15> ), .Y(n184) );
  AOI22X1 U190 ( .A(n182), .B(\w0<15> ), .C(\w1<15> ), .D(n94), .Y(n183) );
endmodule


module four_bank_mem ( clk, rst, createdump, .addr({\addr<15> , \addr<14> , 
        \addr<13> , \addr<12> , \addr<11> , \addr<10> , \addr<9> , \addr<8> , 
        \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> , 
        \addr<1> , \addr<0> }), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        wr, rd, .data_out({\data_out<15> , \data_out<14> , \data_out<13> , 
        \data_out<12> , \data_out<11> , \data_out<10> , \data_out<9> , 
        \data_out<8> , \data_out<7> , \data_out<6> , \data_out<5> , 
        \data_out<4> , \data_out<3> , \data_out<2> , \data_out<1> , 
        \data_out<0> }), stall, .busy({\busy<3> , \busy<2> , \busy<1> , 
        \busy<0> }), err );
  input clk, rst, createdump, \addr<15> , \addr<14> , \addr<13> , \addr<12> ,
         \addr<11> , \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> ,
         \addr<5> , \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> ,
         \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , wr, rd;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , stall,
         \busy<3> , \busy<2> , \busy<1> , \busy<0> , err;
  wire   n109, \en<3> , \en<2> , \en<1> , \en<0> , \data0_out<15> ,
         \data0_out<14> , \data0_out<13> , \data0_out<12> , \data0_out<11> ,
         \data0_out<10> , \data0_out<9> , \data0_out<8> , \data0_out<7> ,
         \data0_out<6> , \data0_out<5> , \data0_out<4> , \data0_out<3> ,
         \data0_out<2> , \data0_out<1> , \data0_out<0> , err0, \data1_out<15> ,
         \data1_out<14> , \data1_out<13> , \data1_out<12> , \data1_out<11> ,
         \data1_out<10> , \data1_out<9> , \data1_out<8> , \data1_out<7> ,
         \data1_out<6> , \data1_out<5> , \data1_out<4> , \data1_out<3> ,
         \data1_out<2> , \data1_out<1> , \data1_out<0> , err1, \data2_out<15> ,
         \data2_out<14> , \data2_out<13> , \data2_out<12> , \data2_out<11> ,
         \data2_out<10> , \data2_out<9> , \data2_out<8> , \data2_out<7> ,
         \data2_out<6> , \data2_out<5> , \data2_out<4> , \data2_out<3> ,
         \data2_out<2> , \data2_out<1> , \data2_out<0> , err2, \data3_out<15> ,
         \data3_out<14> , \data3_out<13> , \data3_out<12> , \data3_out<11> ,
         \data3_out<10> , \data3_out<9> , \data3_out<8> , \data3_out<7> ,
         \data3_out<6> , \data3_out<5> , \data3_out<4> , \data3_out<3> ,
         \data3_out<2> , \data3_out<1> , \data3_out<0> , err3, \bsy0<3> ,
         \bsy0<2> , \bsy0<1> , \bsy0<0> , \bsy1<3> , \bsy1<2> , \bsy1<1> ,
         \bsy1<0> , \bsy2<3> , \bsy2<2> , \bsy2<1> , \bsy2<0> , n8, n9, n10,
         n11, n13, n16, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n1, n2, n3, n4, n5, n6,
         n7, n14, n17, n19, n55, n57, n59, n61, n63, n65, n67, n69, n71, n73,
         n75, n77, n79, n80, n81, n82, n83, n84, n85, n86, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n107, n108;

  NOR3X1 U9 ( .A(n90), .B(n91), .C(n88), .Y(stall) );
  AOI22X1 U10 ( .A(n9), .B(n107), .C(\addr<2> ), .D(n10), .Y(n8) );
  OAI21X1 U11 ( .A(\addr<1> ), .B(n11), .C(n4), .Y(n10) );
  OAI21X1 U13 ( .A(\addr<1> ), .B(n13), .C(n2), .Y(n9) );
  AOI21X1 U15 ( .A(n6), .B(n16), .C(n90), .Y(n109) );
  NOR3X1 U16 ( .A(err1), .B(err3), .C(err2), .Y(n16) );
  NOR3X1 U18 ( .A(n86), .B(\busy<3> ), .C(n90), .Y(\en<3> ) );
  NOR3X1 U20 ( .A(n84), .B(n90), .C(n107), .Y(\en<2> ) );
  NOR3X1 U22 ( .A(n82), .B(n90), .C(n108), .Y(\en<1> ) );
  NOR3X1 U24 ( .A(n80), .B(\busy<0> ), .C(n90), .Y(\en<0> ) );
  NOR2X1 U28 ( .A(\data3_out<9> ), .B(\data2_out<9> ), .Y(n23) );
  NOR2X1 U29 ( .A(\data1_out<9> ), .B(\data0_out<9> ), .Y(n22) );
  NOR2X1 U31 ( .A(\data3_out<8> ), .B(\data2_out<8> ), .Y(n25) );
  NOR2X1 U32 ( .A(\data1_out<8> ), .B(\data0_out<8> ), .Y(n24) );
  NOR2X1 U34 ( .A(\data3_out<7> ), .B(\data2_out<7> ), .Y(n27) );
  NOR2X1 U35 ( .A(\data1_out<7> ), .B(\data0_out<7> ), .Y(n26) );
  NOR2X1 U37 ( .A(\data3_out<6> ), .B(\data2_out<6> ), .Y(n29) );
  NOR2X1 U38 ( .A(\data1_out<6> ), .B(\data0_out<6> ), .Y(n28) );
  NOR2X1 U40 ( .A(\data3_out<5> ), .B(\data2_out<5> ), .Y(n31) );
  NOR2X1 U41 ( .A(\data1_out<5> ), .B(\data0_out<5> ), .Y(n30) );
  NOR2X1 U43 ( .A(\data3_out<4> ), .B(\data2_out<4> ), .Y(n33) );
  NOR2X1 U44 ( .A(\data1_out<4> ), .B(\data0_out<4> ), .Y(n32) );
  NOR2X1 U46 ( .A(\data3_out<3> ), .B(\data2_out<3> ), .Y(n35) );
  NOR2X1 U47 ( .A(\data1_out<3> ), .B(\data0_out<3> ), .Y(n34) );
  NOR2X1 U49 ( .A(\data3_out<2> ), .B(\data2_out<2> ), .Y(n37) );
  NOR2X1 U50 ( .A(\data1_out<2> ), .B(\data0_out<2> ), .Y(n36) );
  NOR2X1 U52 ( .A(\data3_out<1> ), .B(\data2_out<1> ), .Y(n39) );
  NOR2X1 U53 ( .A(\data1_out<1> ), .B(\data0_out<1> ), .Y(n38) );
  NOR2X1 U55 ( .A(\data3_out<15> ), .B(\data2_out<15> ), .Y(n41) );
  NOR2X1 U56 ( .A(\data1_out<15> ), .B(\data0_out<15> ), .Y(n40) );
  NOR2X1 U58 ( .A(\data3_out<14> ), .B(\data2_out<14> ), .Y(n43) );
  NOR2X1 U59 ( .A(\data1_out<14> ), .B(\data0_out<14> ), .Y(n42) );
  NOR2X1 U61 ( .A(\data3_out<13> ), .B(\data2_out<13> ), .Y(n45) );
  NOR2X1 U62 ( .A(\data1_out<13> ), .B(\data0_out<13> ), .Y(n44) );
  NOR2X1 U64 ( .A(\data3_out<12> ), .B(\data2_out<12> ), .Y(n47) );
  NOR2X1 U65 ( .A(\data1_out<12> ), .B(\data0_out<12> ), .Y(n46) );
  NOR2X1 U67 ( .A(\data3_out<11> ), .B(\data2_out<11> ), .Y(n49) );
  NOR2X1 U68 ( .A(\data1_out<11> ), .B(\data0_out<11> ), .Y(n48) );
  NOR2X1 U70 ( .A(\data3_out<10> ), .B(\data2_out<10> ), .Y(n51) );
  NOR2X1 U71 ( .A(\data1_out<10> ), .B(\data0_out<10> ), .Y(n50) );
  NOR2X1 U73 ( .A(\data3_out<0> ), .B(\data2_out<0> ), .Y(n53) );
  NOR2X1 U74 ( .A(\data1_out<0> ), .B(\data0_out<0> ), .Y(n52) );
  NOR3X1 U75 ( .A(\bsy0<3> ), .B(\bsy2<3> ), .C(\bsy1<3> ), .Y(n54) );
  NOR3X1 U76 ( .A(\bsy0<2> ), .B(\bsy2<2> ), .C(\bsy1<2> ), .Y(n11) );
  NOR3X1 U77 ( .A(\bsy0<1> ), .B(\bsy2<1> ), .C(\bsy1<1> ), .Y(n20) );
  NOR3X1 U78 ( .A(\bsy0<0> ), .B(\bsy2<0> ), .C(\bsy1<0> ), .Y(n13) );
  final_memory_3 m0 ( .data_out({\data0_out<15> , \data0_out<14> , 
        \data0_out<13> , \data0_out<12> , \data0_out<11> , \data0_out<10> , 
        \data0_out<9> , \data0_out<8> , \data0_out<7> , \data0_out<6> , 
        \data0_out<5> , \data0_out<4> , \data0_out<3> , \data0_out<2> , 
        \data0_out<1> , \data0_out<0> }), .err(err0), .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<15> , \addr<14> , \addr<13> , \addr<12> , 
        \addr<11> , \addr<10> , \addr<9> , \addr<8> , n101, n99, n97, n95, n93}), .wr(wr), .rd(rd), .enable(\en<0> ), .create_dump(createdump), .bank_id({
        1'b0, 1'b0}), .clk(clk), .rst(n91) );
  final_memory_2 m1 ( .data_out({\data1_out<15> , \data1_out<14> , 
        \data1_out<13> , \data1_out<12> , \data1_out<11> , \data1_out<10> , 
        \data1_out<9> , \data1_out<8> , \data1_out<7> , \data1_out<6> , 
        \data1_out<5> , \data1_out<4> , \data1_out<3> , \data1_out<2> , 
        \data1_out<1> , \data1_out<0> }), .err(err1), .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<15> , \addr<14> , \addr<13> , \addr<12> , 
        \addr<11> , \addr<10> , \addr<9> , \addr<8> , n101, n99, n97, n95, n93}), .wr(wr), .rd(rd), .enable(\en<1> ), .create_dump(createdump), .bank_id({
        1'b0, 1'b1}), .clk(clk), .rst(n91) );
  final_memory_1 m2 ( .data_out({\data2_out<15> , \data2_out<14> , 
        \data2_out<13> , \data2_out<12> , \data2_out<11> , \data2_out<10> , 
        \data2_out<9> , \data2_out<8> , \data2_out<7> , \data2_out<6> , 
        \data2_out<5> , \data2_out<4> , \data2_out<3> , \data2_out<2> , 
        \data2_out<1> , \data2_out<0> }), .err(err2), .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<15> , \addr<14> , \addr<13> , \addr<12> , 
        \addr<11> , \addr<10> , \addr<9> , \addr<8> , n101, n99, n97, n95, n93}), .wr(wr), .rd(rd), .enable(\en<2> ), .create_dump(createdump), .bank_id({
        1'b1, 1'b0}), .clk(clk), .rst(n91) );
  final_memory_0 m3 ( .data_out({\data3_out<15> , \data3_out<14> , 
        \data3_out<13> , \data3_out<12> , \data3_out<11> , \data3_out<10> , 
        \data3_out<9> , \data3_out<8> , \data3_out<7> , \data3_out<6> , 
        \data3_out<5> , \data3_out<4> , \data3_out<3> , \data3_out<2> , 
        \data3_out<1> , \data3_out<0> }), .err(err3), .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<15> , \addr<14> , \addr<13> , \addr<12> , 
        \addr<11> , \addr<10> , \addr<9> , \addr<8> , n101, n99, n97, n95, n93}), .wr(wr), .rd(rd), .enable(\en<3> ), .create_dump(createdump), .bank_id({
        1'b1, 1'b1}), .clk(clk), .rst(n91) );
  dff_216 \b0[0]  ( .q(\bsy0<0> ), .d(\en<0> ), .clk(clk), .rst(n91) );
  dff_217 \b0[1]  ( .q(\bsy0<1> ), .d(\en<1> ), .clk(clk), .rst(n91) );
  dff_218 \b0[2]  ( .q(\bsy0<2> ), .d(\en<2> ), .clk(clk), .rst(n91) );
  dff_219 \b0[3]  ( .q(\bsy0<3> ), .d(\en<3> ), .clk(clk), .rst(n91) );
  dff_212 \b1[0]  ( .q(\bsy1<0> ), .d(\bsy0<0> ), .clk(clk), .rst(n91) );
  dff_213 \b1[1]  ( .q(\bsy1<1> ), .d(\bsy0<1> ), .clk(clk), .rst(n91) );
  dff_214 \b1[2]  ( .q(\bsy1<2> ), .d(\bsy0<2> ), .clk(clk), .rst(n91) );
  dff_215 \b1[3]  ( .q(\bsy1<3> ), .d(\bsy0<3> ), .clk(clk), .rst(n91) );
  dff_208 \b2[0]  ( .q(\bsy2<0> ), .d(\bsy1<0> ), .clk(clk), .rst(n91) );
  dff_209 \b2[1]  ( .q(\bsy2<1> ), .d(\bsy1<1> ), .clk(clk), .rst(n91) );
  dff_210 \b2[2]  ( .q(\bsy2<2> ), .d(\bsy1<2> ), .clk(clk), .rst(n91) );
  dff_211 \b2[3]  ( .q(\bsy2<3> ), .d(\bsy1<3> ), .clk(clk), .rst(n91) );
  INVX1 U3 ( .A(rst), .Y(n92) );
  INVX1 U4 ( .A(n54), .Y(\busy<3> ) );
  OR2X1 U5 ( .A(err0), .B(\addr<0> ), .Y(n5) );
  INVX1 U6 ( .A(n94), .Y(n93) );
  INVX1 U7 ( .A(n96), .Y(n95) );
  INVX1 U8 ( .A(n98), .Y(n97) );
  INVX1 U12 ( .A(n100), .Y(n99) );
  INVX1 U14 ( .A(\addr<6> ), .Y(n100) );
  INVX1 U17 ( .A(n102), .Y(n101) );
  INVX1 U19 ( .A(\addr<7> ), .Y(n102) );
  INVX1 U21 ( .A(\addr<1> ), .Y(n108) );
  INVX1 U23 ( .A(\addr<2> ), .Y(n107) );
  INVX1 U25 ( .A(n20), .Y(\busy<1> ) );
  INVX1 U26 ( .A(n13), .Y(\busy<0> ) );
  INVX1 U27 ( .A(n11), .Y(\busy<2> ) );
  INVX1 U30 ( .A(\addr<5> ), .Y(n98) );
  INVX1 U33 ( .A(n92), .Y(n91) );
  AND2X1 U36 ( .A(\addr<1> ), .B(\busy<1> ), .Y(n1) );
  INVX1 U39 ( .A(n1), .Y(n2) );
  AND2X1 U42 ( .A(\addr<1> ), .B(\busy<3> ), .Y(n3) );
  INVX1 U45 ( .A(n3), .Y(n4) );
  INVX1 U48 ( .A(n5), .Y(n6) );
  AND2X2 U51 ( .A(n52), .B(n53), .Y(n7) );
  INVX1 U54 ( .A(n7), .Y(\data_out<0> ) );
  AND2X2 U57 ( .A(n50), .B(n51), .Y(n14) );
  INVX1 U60 ( .A(n14), .Y(\data_out<10> ) );
  AND2X2 U63 ( .A(n48), .B(n49), .Y(n17) );
  INVX1 U66 ( .A(n17), .Y(\data_out<11> ) );
  AND2X2 U69 ( .A(n46), .B(n47), .Y(n19) );
  INVX1 U72 ( .A(n19), .Y(\data_out<12> ) );
  AND2X2 U79 ( .A(n44), .B(n45), .Y(n55) );
  INVX1 U80 ( .A(n55), .Y(\data_out<13> ) );
  AND2X2 U81 ( .A(n42), .B(n43), .Y(n57) );
  INVX1 U82 ( .A(n57), .Y(\data_out<14> ) );
  AND2X2 U83 ( .A(n40), .B(n41), .Y(n59) );
  INVX1 U84 ( .A(n59), .Y(\data_out<15> ) );
  AND2X2 U85 ( .A(n38), .B(n39), .Y(n61) );
  INVX1 U86 ( .A(n61), .Y(\data_out<1> ) );
  AND2X2 U87 ( .A(n36), .B(n37), .Y(n63) );
  INVX1 U88 ( .A(n63), .Y(\data_out<2> ) );
  AND2X2 U89 ( .A(n34), .B(n35), .Y(n65) );
  INVX1 U90 ( .A(n65), .Y(\data_out<3> ) );
  AND2X2 U91 ( .A(n32), .B(n33), .Y(n67) );
  INVX1 U92 ( .A(n67), .Y(\data_out<4> ) );
  AND2X2 U93 ( .A(n30), .B(n31), .Y(n69) );
  INVX1 U94 ( .A(n69), .Y(\data_out<5> ) );
  AND2X2 U95 ( .A(n28), .B(n29), .Y(n71) );
  INVX1 U96 ( .A(n71), .Y(\data_out<6> ) );
  AND2X2 U97 ( .A(n26), .B(n27), .Y(n73) );
  INVX1 U98 ( .A(n73), .Y(\data_out<7> ) );
  AND2X2 U99 ( .A(n24), .B(n25), .Y(n75) );
  INVX1 U100 ( .A(n75), .Y(\data_out<8> ) );
  AND2X2 U101 ( .A(n22), .B(n23), .Y(n77) );
  INVX1 U102 ( .A(n77), .Y(\data_out<9> ) );
  AND2X1 U103 ( .A(n108), .B(n107), .Y(n79) );
  INVX1 U104 ( .A(n79), .Y(n80) );
  AND2X1 U105 ( .A(n20), .B(n107), .Y(n81) );
  INVX1 U106 ( .A(n81), .Y(n82) );
  AND2X1 U107 ( .A(n11), .B(n108), .Y(n83) );
  INVX1 U108 ( .A(n83), .Y(n84) );
  AND2X1 U109 ( .A(\addr<2> ), .B(\addr<1> ), .Y(n85) );
  INVX1 U110 ( .A(n85), .Y(n86) );
  BUFX2 U111 ( .A(n109), .Y(err) );
  BUFX2 U112 ( .A(n8), .Y(n88) );
  OR2X1 U113 ( .A(rd), .B(wr), .Y(n89) );
  INVX1 U114 ( .A(n89), .Y(n90) );
  INVX1 U115 ( .A(\addr<4> ), .Y(n96) );
  INVX1 U116 ( .A(\addr<3> ), .Y(n94) );
endmodule


module mem_system_control ( clk, rst, rd, wr, hit, dirty, cache_wr, cache_hit, 
        cache_sel, .cache_offset({\cache_offset<1> , \cache_offset<0> }), comp, 
        stall, err, done, mem_rd, mem_wr, mem_sel, .mem_offset({
        \mem_offset<1> , \mem_offset<0> }) );
  input clk, rst, rd, wr, hit, dirty;
  output cache_wr, cache_hit, cache_sel, \cache_offset<1> , \cache_offset<0> ,
         comp, stall, err, done, mem_rd, mem_wr, mem_sel, \mem_offset<1> ,
         \mem_offset<0> ;


  mem_state_reg STATE_FF ( .clk(clk), .rst(rst), .state({1'b0, 1'b0, 1'b0, 
        1'b0}), .next_state() );
  mem_next_state NEXT_STATE ( .rd(rd), .wr(wr), .hit(hit), .dirty(dirty), 
        .state({1'b0, 1'b0, 1'b0, 1'b0}), .err(err), .next_state() );
  mem_signals SIGNALS ( .hit(hit), .state({1'b0, 1'b0, 1'b0, 1'b0}), .stall(
        stall), .done(done), .cache_wr(cache_wr), .cache_hit(cache_hit), 
        .cache_offset({\cache_offset<1> , \cache_offset<0> }), .cache_sel(
        cache_sel), .comp(comp), .mem_wr(mem_wr), .mem_rd(mem_rd), 
        .mem_offset({\mem_offset<1> , \mem_offset<0> }), .mem_sel(mem_sel) );
endmodule


module mem_system ( .DataOut({\DataOut<15> , \DataOut<14> , \DataOut<13> , 
        \DataOut<12> , \DataOut<11> , \DataOut<10> , \DataOut<9> , 
        \DataOut<8> , \DataOut<7> , \DataOut<6> , \DataOut<5> , \DataOut<4> , 
        \DataOut<3> , \DataOut<2> , \DataOut<1> , \DataOut<0> }), Done, Stall, 
        CacheHit, err, .Addr({\Addr<15> , \Addr<14> , \Addr<13> , \Addr<12> , 
        \Addr<11> , \Addr<10> , \Addr<9> , \Addr<8> , \Addr<7> , \Addr<6> , 
        \Addr<5> , \Addr<4> , \Addr<3> , \Addr<2> , \Addr<1> , \Addr<0> }), 
    .DataIn({\DataIn<15> , \DataIn<14> , \DataIn<13> , \DataIn<12> , 
        \DataIn<11> , \DataIn<10> , \DataIn<9> , \DataIn<8> , \DataIn<7> , 
        \DataIn<6> , \DataIn<5> , \DataIn<4> , \DataIn<3> , \DataIn<2> , 
        \DataIn<1> , \DataIn<0> }), Rd, Wr, createdump, clk, rst );
  input \Addr<15> , \Addr<14> , \Addr<13> , \Addr<12> , \Addr<11> , \Addr<10> ,
         \Addr<9> , \Addr<8> , \Addr<7> , \Addr<6> , \Addr<5> , \Addr<4> ,
         \Addr<3> , \Addr<2> , \Addr<1> , \Addr<0> , \DataIn<15> ,
         \DataIn<14> , \DataIn<13> , \DataIn<12> , \DataIn<11> , \DataIn<10> ,
         \DataIn<9> , \DataIn<8> , \DataIn<7> , \DataIn<6> , \DataIn<5> ,
         \DataIn<4> , \DataIn<3> , \DataIn<2> , \DataIn<1> , \DataIn<0> , Rd,
         Wr, createdump, clk, rst;
  output \DataOut<15> , \DataOut<14> , \DataOut<13> , \DataOut<12> ,
         \DataOut<11> , \DataOut<10> , \DataOut<9> , \DataOut<8> ,
         \DataOut<7> , \DataOut<6> , \DataOut<5> , \DataOut<4> , \DataOut<3> ,
         \DataOut<2> , \DataOut<1> , \DataOut<0> , Done, Stall, CacheHit, err;
  wire   cache_sel, cache_write, cache_wr, \mem_data_out<15> ,
         \mem_data_out<14> , \mem_data_out<13> , \mem_data_out<12> ,
         \mem_data_out<11> , \mem_data_out<10> , \mem_data_out<9> ,
         \mem_data_out<8> , \mem_data_out<7> , \mem_data_out<6> ,
         \mem_data_out<5> , \mem_data_out<4> , \mem_data_out<3> ,
         \mem_data_out<2> , \mem_data_out<1> , \mem_data_out<0> ,
         \cache_offset<1> , \cache_offset<0> , \cache_off<0> , mem_sel,
         mem_addr_2, mem_addr_1, \cache_tag_out<4> , \cache_tag_out<3> ,
         \cache_tag_out<2> , \cache_tag_out<1> , \cache_tag_out<0> , cache_hit,
         cache_dirty, cache_valid, cache_err, _0_net_, comp, mem_err, mem_wr,
         mem_rd, control_err, _2_net_, n29, n30, n31, n32, n33, n34, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120;

  OR2X2 U5 ( .A(Rd), .B(Wr), .Y(_0_net_) );
  AOI22X1 U33 ( .A(mem_sel), .B(\Addr<15> ), .C(\cache_tag_out<4> ), .D(n119), 
        .Y(n29) );
  AOI22X1 U34 ( .A(\Addr<14> ), .B(mem_sel), .C(\cache_tag_out<3> ), .D(n119), 
        .Y(n30) );
  AOI22X1 U35 ( .A(\Addr<13> ), .B(mem_sel), .C(\cache_tag_out<2> ), .D(n119), 
        .Y(n31) );
  AOI22X1 U36 ( .A(\Addr<12> ), .B(mem_sel), .C(\cache_tag_out<1> ), .D(n119), 
        .Y(n32) );
  AOI22X1 U37 ( .A(\Addr<11> ), .B(mem_sel), .C(\cache_tag_out<0> ), .D(n119), 
        .Y(n33) );
  NOR3X1 U38 ( .A(cache_err), .B(mem_err), .C(control_err), .Y(n34) );
  OAI21X1 U39 ( .A(n84), .B(n120), .C(n57), .Y(cache_write) );
  AOI22X1 U41 ( .A(\Addr<2> ), .B(n118), .C(\cache_offset<1> ), .D(n83), .Y(
        n36) );
  AOI22X1 U42 ( .A(\Addr<1> ), .B(n118), .C(\cache_offset<0> ), .D(n83), .Y(
        n37) );
  AOI22X1 U43 ( .A(\DataIn<9> ), .B(n118), .C(\mem_data_out<9> ), .D(n83), .Y(
        n38) );
  AOI22X1 U44 ( .A(\DataIn<8> ), .B(n118), .C(\mem_data_out<8> ), .D(n83), .Y(
        n39) );
  AOI22X1 U45 ( .A(\DataIn<7> ), .B(n118), .C(\mem_data_out<7> ), .D(n83), .Y(
        n40) );
  AOI22X1 U46 ( .A(\DataIn<6> ), .B(n118), .C(\mem_data_out<6> ), .D(n83), .Y(
        n41) );
  AOI22X1 U47 ( .A(\DataIn<5> ), .B(n118), .C(\mem_data_out<5> ), .D(n83), .Y(
        n42) );
  AOI22X1 U48 ( .A(\DataIn<4> ), .B(n118), .C(\mem_data_out<4> ), .D(n83), .Y(
        n43) );
  AOI22X1 U49 ( .A(\DataIn<3> ), .B(n118), .C(\mem_data_out<3> ), .D(n84), .Y(
        n44) );
  AOI22X1 U50 ( .A(\DataIn<2> ), .B(n118), .C(\mem_data_out<2> ), .D(n84), .Y(
        n45) );
  AOI22X1 U51 ( .A(\DataIn<1> ), .B(n118), .C(\mem_data_out<1> ), .D(n84), .Y(
        n46) );
  AOI22X1 U52 ( .A(\DataIn<15> ), .B(n118), .C(\mem_data_out<15> ), .D(n84), 
        .Y(n47) );
  AOI22X1 U53 ( .A(\DataIn<14> ), .B(n118), .C(\mem_data_out<14> ), .D(n84), 
        .Y(n48) );
  AOI22X1 U54 ( .A(\DataIn<13> ), .B(n118), .C(\mem_data_out<13> ), .D(n84), 
        .Y(n49) );
  AOI22X1 U55 ( .A(\DataIn<12> ), .B(n118), .C(\mem_data_out<12> ), .D(n84), 
        .Y(n50) );
  AOI22X1 U56 ( .A(\DataIn<11> ), .B(n118), .C(\mem_data_out<11> ), .D(n84), 
        .Y(n51) );
  AOI22X1 U57 ( .A(\DataIn<10> ), .B(n118), .C(\mem_data_out<10> ), .D(n84), 
        .Y(n52) );
  AOI22X1 U58 ( .A(\DataIn<0> ), .B(n118), .C(\mem_data_out<0> ), .D(n84), .Y(
        n53) );
  cache_cache_id0 c0 ( .enable(_0_net_), .clk(clk), .rst(n85), .createdump(
        createdump), .tag_in({\Addr<15> , \Addr<14> , \Addr<13> , \Addr<12> , 
        \Addr<11> }), .index({n82, n81, n80, n92, n90, n88, \Addr<4> , n79}), 
        .offset({n116, n117, \cache_off<0> }), .data_in({n110, n109, n108, 
        n107, n106, n105, n104, n103, n102, n101, n100, n99, n98, n97, n96, 
        n95}), .comp(comp), .write(cache_write), .valid_in(1'b1), .tag_out({
        \cache_tag_out<4> , \cache_tag_out<3> , \cache_tag_out<2> , 
        \cache_tag_out<1> , \cache_tag_out<0> }), .data_out({\DataOut<15> , 
        \DataOut<14> , \DataOut<13> , \DataOut<12> , \DataOut<11> , 
        \DataOut<10> , \DataOut<9> , \DataOut<8> , \DataOut<7> , \DataOut<6> , 
        \DataOut<5> , \DataOut<4> , \DataOut<3> , \DataOut<2> , \DataOut<1> , 
        \DataOut<0> }), .hit(cache_hit), .dirty(cache_dirty), .valid(
        cache_valid), .err(cache_err) );
  four_bank_mem mem ( .clk(clk), .rst(n85), .createdump(createdump), .addr({
        n111, n112, n113, n114, n115, n82, n81, n80, n92, n90, n88, n55, n54, 
        mem_addr_2, mem_addr_1, 1'b0}), .data_in({\DataOut<15> , \DataOut<14> , 
        \DataOut<13> , \DataOut<12> , \DataOut<11> , \DataOut<10> , 
        \DataOut<9> , \DataOut<8> , \DataOut<7> , \DataOut<6> , \DataOut<5> , 
        \DataOut<4> , \DataOut<3> , \DataOut<2> , \DataOut<1> , \DataOut<0> }), 
        .wr(mem_wr), .rd(mem_rd), .data_out({\mem_data_out<15> , 
        \mem_data_out<14> , \mem_data_out<13> , \mem_data_out<12> , 
        \mem_data_out<11> , \mem_data_out<10> , \mem_data_out<9> , 
        \mem_data_out<8> , \mem_data_out<7> , \mem_data_out<6> , 
        \mem_data_out<5> , \mem_data_out<4> , \mem_data_out<3> , 
        \mem_data_out<2> , \mem_data_out<1> , \mem_data_out<0> }), .stall(), 
        .busy(), .err(mem_err) );
  mem_system_control ctl ( .clk(clk), .rst(n85), .rd(Rd), .wr(Wr), .hit(
        _2_net_), .dirty(cache_dirty), .cache_wr(cache_wr), .cache_hit(
        CacheHit), .cache_sel(cache_sel), .cache_offset({\cache_offset<1> , 
        \cache_offset<0> }), .comp(comp), .stall(Stall), .err(control_err), 
        .done(Done), .mem_rd(mem_rd), .mem_wr(mem_wr), .mem_sel(mem_sel), 
        .mem_offset({mem_addr_2, mem_addr_1}) );
  INVX1 U59 ( .A(Wr), .Y(n120) );
  AND2X1 U60 ( .A(\Addr<0> ), .B(n118), .Y(\cache_off<0> ) );
  BUFX2 U61 ( .A(\Addr<8> ), .Y(n80) );
  BUFX2 U62 ( .A(\Addr<10> ), .Y(n82) );
  BUFX2 U63 ( .A(cache_sel), .Y(n84) );
  BUFX2 U64 ( .A(cache_sel), .Y(n83) );
  INVX1 U65 ( .A(n83), .Y(n118) );
  INVX1 U66 ( .A(\Addr<5> ), .Y(n89) );
  INVX1 U67 ( .A(\Addr<6> ), .Y(n91) );
  INVX1 U68 ( .A(\Addr<7> ), .Y(n93) );
  INVX1 U69 ( .A(mem_sel), .Y(n119) );
  AND2X1 U70 ( .A(cache_valid), .B(cache_hit), .Y(_2_net_) );
  INVX1 U71 ( .A(n34), .Y(err) );
  INVX1 U72 ( .A(n89), .Y(n88) );
  BUFX2 U73 ( .A(n79), .Y(n54) );
  BUFX2 U74 ( .A(\Addr<4> ), .Y(n55) );
  INVX2 U75 ( .A(rst), .Y(n86) );
  INVX8 U76 ( .A(n87), .Y(n79) );
  INVX2 U77 ( .A(\Addr<3> ), .Y(n87) );
  AND2X1 U78 ( .A(cache_wr), .B(n84), .Y(n56) );
  INVX1 U79 ( .A(n56), .Y(n57) );
  BUFX2 U80 ( .A(n53), .Y(n58) );
  INVX1 U81 ( .A(n58), .Y(n95) );
  BUFX2 U82 ( .A(n52), .Y(n59) );
  INVX1 U83 ( .A(n59), .Y(n105) );
  BUFX2 U84 ( .A(n51), .Y(n60) );
  INVX1 U85 ( .A(n60), .Y(n106) );
  BUFX2 U86 ( .A(n50), .Y(n61) );
  INVX1 U87 ( .A(n61), .Y(n107) );
  BUFX2 U88 ( .A(n49), .Y(n62) );
  INVX1 U89 ( .A(n62), .Y(n108) );
  BUFX2 U90 ( .A(n48), .Y(n63) );
  INVX1 U91 ( .A(n63), .Y(n109) );
  BUFX2 U92 ( .A(n47), .Y(n64) );
  INVX1 U93 ( .A(n64), .Y(n110) );
  BUFX2 U94 ( .A(n46), .Y(n65) );
  INVX1 U95 ( .A(n65), .Y(n96) );
  BUFX2 U96 ( .A(n45), .Y(n66) );
  INVX1 U97 ( .A(n66), .Y(n97) );
  BUFX2 U98 ( .A(n44), .Y(n67) );
  INVX1 U99 ( .A(n67), .Y(n98) );
  BUFX2 U100 ( .A(n43), .Y(n68) );
  INVX1 U101 ( .A(n68), .Y(n99) );
  BUFX2 U102 ( .A(n42), .Y(n69) );
  INVX1 U103 ( .A(n69), .Y(n100) );
  BUFX2 U104 ( .A(n41), .Y(n70) );
  INVX1 U105 ( .A(n70), .Y(n101) );
  BUFX2 U106 ( .A(n40), .Y(n71) );
  INVX1 U107 ( .A(n71), .Y(n102) );
  BUFX2 U108 ( .A(n39), .Y(n72) );
  INVX1 U109 ( .A(n72), .Y(n103) );
  BUFX2 U110 ( .A(n38), .Y(n73) );
  INVX1 U111 ( .A(n73), .Y(n104) );
  BUFX2 U112 ( .A(n36), .Y(n74) );
  INVX1 U113 ( .A(n74), .Y(n116) );
  BUFX2 U114 ( .A(n33), .Y(n75) );
  INVX1 U115 ( .A(n75), .Y(n115) );
  BUFX2 U116 ( .A(n32), .Y(n76) );
  INVX1 U117 ( .A(n76), .Y(n114) );
  INVX1 U118 ( .A(n31), .Y(n113) );
  BUFX2 U119 ( .A(n30), .Y(n77) );
  INVX1 U120 ( .A(n77), .Y(n112) );
  BUFX2 U121 ( .A(n29), .Y(n78) );
  INVX1 U122 ( .A(n78), .Y(n111) );
  BUFX2 U123 ( .A(\Addr<9> ), .Y(n81) );
  INVX1 U124 ( .A(n37), .Y(n117) );
  INVX8 U125 ( .A(n86), .Y(n85) );
  INVX8 U126 ( .A(n91), .Y(n90) );
  INVX8 U127 ( .A(n93), .Y(n92) );
endmodule

