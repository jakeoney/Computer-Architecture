library verilog;
use verilog.vl_types.all;
entity shifter_hier_bench is
end shifter_hier_bench;
